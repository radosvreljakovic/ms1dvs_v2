// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tCAaz71uuf6m2PfNJraOUwRM/qHIPOu7nO9Rbj6DvaZ7VbfP6A5MKZRg4YgDYNIr
SD0DZRMECvgZkTnciyj9pPIozr5d7tYVa2OdHw4hGzhswvgJEI+KUzr72uWAS3UT
AxUwR5fJhdCnzuIAQLp1ljKRMZTdJtQKpT2N+iL/tl4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13472)
gDR9cKjn3XSrwGhP00hhNJYMc+0syEB9wBP/Cmh/S7wnazK4CRPlNSyjpyKrmdML
8+2wCuLzveCcQBHqHGzoW+nhh519zYv16s2xBMRhaZdZc6ez6iXi1+MFADOagoQj
eyu6NWJxQIlRSL/dVO+HBknTeyefVzN9W3V3AuCe7MpIDs2YsLw2iqAGlJNzIz73
8hM7q0wsUMK5aj4CE4tTObKnbEVrLqv7abWzRmGog87+M9qgxKcWC2jxn607ant4
5QjNsO05STyINqfwEodEYCJ40ZXBy/i5GEDN7c8LHLRcvxe7l8jcsSkiNpFTBFho
mnuyNx0dA4FDPvCHrGZ4YGD1pynGswDV6dNxBZJOoa2UYR06qbv0oh2ykuPM7SW8
6o4e0x+jvpbCTXLhdHYFzCIRoT8QPn7OT8t+5EDYNPAMSoWLq/yQAykwLO55BBdR
YDRHrJ9RQVavtXThpCWt1t8b0tqra7ZzqyTgvcsX4/v1WnAv5TiJn5VgwavY+4aa
yM31m809LnyZhAoJdN9q1uWll9WctfQXjCcFh+mCVQY15Vb3pKUDT+BBZfOTi9qV
UJwXsMnzOM2XHcaTuGxzZ8V2ZhZCgw5B+UsGfhs0RGk3Ye56RtGAH/nA7Y+hiVi0
ZmSA/8sWTg4jK+FxuQ5IrH4LlRgIKJT5CSqh57jYb3c87PtEsHCFzejkZ8DPdsS9
feUHQ5/Qx0se+w3O5adN4HBAAG0agnYLSWqNSZu+UR0DhWJFZYMLARnS2CiObOtI
aiJvQ840BfXore3EFsE6ry7zvuZTLQvLlSZkDYYMSj8cOUZGwkem7bHRgovd8tF4
Iec3h7do5Wfflp9IXJEeU5edW+Mp5WvAEiB7ySg9GDAEq0W6EFCt1MT3gvMANGJI
M13ExvKzDWdBIbVsZ7W8cKv4QTtlbx0DZxph//Qbkw4pmR/CphidJoUDWqTwF3t6
3x2a7AUD37hkTnBhPyMXmqdRNOZPrKCoTuLUZi/thiFrQv5FDwd8wfte1d2QqvYa
ApG9c4ORJwGj6XShzeBsWP5Qi+foP5Qt/mRNGifrW6DaYiVwVGgv1i2f1XsNRrkg
debd6Q82JtSDSpLEs2dxsBHD5LbdpuAghpktvEEeg9M+Mf4/o8yatsZlVq8cns33
ZqzspfVadL6/veYuaqmHvOKFOAnsuC6NfK6S6xLhBJq7mHDgf9hUolhCqHuWl/FD
DEWsCLGI8I7yKXWUeWsb/hnR8Jtveppf8bmYYRZluI3WbZD9SIrH7XLXeeVCwbzc
6MlsUTK+rk/nZIp4YNaiLdbnwe5/cxsHlk5J64BhLY3Ga3AtqgNxW91hvY2loKOs
8pP3HDj8w150Sn1XNFfmgAq7p/QqfOXgjpqauUqjglTutsouMj/VHfkSFI/kjY8p
44wDr2B0Qu0cX+obe8MIVzFT1bmRjxj/XeSi6cmIjCqSFTJHEGZPdq3yAAkdaySA
mxv8sYYB2cVV+yOIWL/eIoXO3S8jm2IbwXH3XqT03V1ZTB0AZ7p0/RnzQXLNflas
YqgM0Du3I00FVnti4/3sMYgAtoFLwzMX9tVFvrd6gsVgrWE0HvmeNe51NDeX8ZUP
d5OBkZpy9AY2R9GhmhFy++uBwDdcDYom4woecwmym3J9z9YwXtHZjCOJvTIgL1WZ
g7FJrwWMSbEY++seTH/tOjgF9Q+e+GkTwDxAkErPHnnBWfwKMGZSTqwFFs+yPRLq
ueYerDwdyf+O8WRf94WCRSpbRp1W6EXu4UPDVMae1veFc5T6Pec9JXy7Zz7PvQ/y
le/bR+K214cEDb9L63W7MT5xTYGlcUgDuCaR6nCNPVGOPsZkYL/Mk2/lwFMkrx0b
wHKxiYYKNpMmV1ICkfZpWVuAqHOYap57Uf6kJ1bNPF+ylRO7CZtvLePuaBEjnb4l
pVYS5NJRtPace1c/URhDFGfegJtTlw54GGnJRMTZJCU8DgSb67cGaZ5kq7XHgruM
uPpXUlCFqXz7hmSOogZfHABOOYClu7FrAiskgQ/6vWMwSUAOFI1wkGXxgPqyKALp
Xq9s24Rkc2s6aBNyOkFle21Xlqpu0B1mv/YJEVjM0ws9nQ0uBcr3sEzzTSUsCank
ZhWYsM3/b9fEfFmaLY80hR+w7B7tW1Uy1oht7+WHsTaGW96RaSY07jENnUF0zbso
9K9DCSMGWfKjutfHHNJtrGx6vFegxwi+2L0LEBSdujeBtoP1os3eATrBqC0bKC+B
L5L5TPc2BSgY0AFY9/o6XU0FnnlddCDAlNQu4G1I6INQ64aGBl+LLiUv1J9FLJfv
ptMQ/OlREdmfhQu+Fy9+eFK5V5JzP88/fUPVAyJcJiqQReG5q3CrLKQrRQhVLs+P
npx53ZCOA4GQ1lVgokLf6JicWmOF/+xNGNHqOvncNYban9w8VWktYPj5+pDZKkmu
2WF8lW5FRiRzcdlHQkWwb2SeECbc3OOmsCeHlknffTqBVumaoW8zbioN2H5BtBim
Il01OwpagZ/hPvQTCWAaEvMQKJY+TY67dfip/N3X6ihjtGG74g+a/5xqgHG6BsvQ
JxL6wyLy7GlYQLMWUYzyX0EGSH3iCiL0/MOwzILVe7snu/KkJI5Wt8EBRzFAorSe
31GVu7olK1dLk2ShN9ZeM2MiBUkR+8HGZxmAk4FG6fUpDCeTpu4J7nrHUuU18nB5
RHmfvRZPQaebJHA8hyA0FTkTLyg/gIlLHcof5bcTbE019hZEqe79Brhk90aDecsw
C93goRyqoJ0WfddRCEELiNnaFbaggIs27qXZhntF9aHa30UrDFD6fxzWR16vR1RA
z9/Wq+8E+hrQVps4Lvo4y+s9JDCQejc6Tmn6iHuLMQDMfQSHDX02TbAFN+SZeuix
InFdaam04dh7aoUKp2vfMs8K37t0GZNMRbz78p8SMIxnd+nCjxjJCzt0Y3IeFm/k
bB6VZR4YKPYOClAH93m94tWF573s5OzpgLR47mHF7BYPTqcuyUgdy4uvMzpxpVI2
52aYu/PuiNjho8Lwv1nDaCo5flZrkQ9KXlBmCGmEds39ZYXsJZQh9pBuKR9k4SMu
hzZo0IJbyvY51cbmtvdNOYx1yms4neb5XFypLMe3QYp8MRgBHR2N87jja9ZXnjx1
T7RNNnuvXqSaTpLIB1Ck8mpEh9mEb0uLfkVhrJbGBO0e/K0ulk94Ow/iY6v5VHJg
4P/JsrMXVA1NO7Dhpxw1EGMvMzb8IWIhaT48sASbpgPozTUSU8XkiF9NTjUz0bst
r/+QxMLU2OEKHsc7Pwtb8jsTIirHQAW7YnlqT0Nni8FXSGIeT6ar0/op/JiHCDU1
ybBo76gMt4q4/6F2oKFaP4vm21bPu8ATsApv8v0DAslSdRxG3JgZsN/0cvUAj/cc
g6/23k2Ohgwz1xCEenokfMrrFCFOGQ4rHFSXzcgLC8jT+nEVIUaOezHwLgkrEH+2
ewhQUb3efgMxE5/zUwV88AeufWL51NVxVN+dV4orfLUteWSbfZSby77Y+E7n8UbK
kpx20bGWCGjyFb3BdVNSf6vste6NSBt9NYIdro1v3NIogU98gS4BpHkd4GApe1k8
/Enj4kjuSRqod0jY6jSigtG94qolkWKYXgYDUgxnSQPYgzQTD8XxUSUCO0D5opFU
oti3G7498QzYmAKVguIZV3rGslxjpzBkmM32cW37i43InNiGpDPYE8p0RPtF79sC
+9UauxBPU0fL9y9oz5U2PKUvvT5BhZ3RlIQMK7hxrvLtp6hh1zar05IWeUjx1CgN
l1XZOXJ3JI4hX+qHOv+sHvgC2CEbLQbEUiK0nWoLR1+OW8LjIpGpPuQWSgx35upk
P3e1ta681+7/ranCrrcYrwyDBZKuILgWBEuK5splP5zHwrI5Bh/4G5mAmehju6On
KssgUvWCXmFkquzKLq6rVNKnI2lR7XElLoVKT+Drhj6xCDnwzi7CiSvz+9dNBi5F
HNaAKFa7yeIeOJhkXRRqYuvNytfYT2xyZkdVAbSU9Oh9T1ctAJo9qilqoB3r4XT5
+0uqTmyUhVuYMbPYPfV5Fp7I02mf0lufqQV9ko4k6nhR+tzu11Stb7PUiS/STXk5
mSj4wZBb8/SD/uoJp89pewQF7CTCbKJglW6a+zDZrGWiSzIZDva1YBSxwlj7QS75
iBy4SjLZ84k2qoVhLhTKT788v9OOhCpYulATINFZl0uGnEOuqZ6IP6qJx2MpLOjX
/Io3o9GLnYAIEzbgGBncXmbUauzVNQyoG/WuzOekaJiFhghGwGt66nrnSXsy6t/M
oJk5cCGY7DCVbnBz1EwuxV5DFHFGd+EdyZE7unRGuSZXD1prYDkPhkxi9N3uVzzl
//if2jwKXfJOMwLwiH+4oHozqJiORnIyb9Q5wqHnDzM8lbayyB/O9TIsVuHY0eB8
ObY+Yp2Lh3jcL8jiP6LJu+dYLrQGd1fd5cwfQ+0z7hNYIaLLP2A7bSl5gsflspU3
9mYtNro7aGlqcETDbXawg24oAtiFl/RX8acO/t1uOeaITfh1SwgVaEJY6fT94M+h
wEnyztGul/M8JT06lfuppOezWgzJpqtKizyMB5l1mTxP70IWpbu3lP6efuGIT1NR
b5R26m1KCxviKYPc2a+GxHNeY/3ZaTacukBwBwQXJaKJLhQvNo8zYR6zUHrUjf6b
aBHPCU1BV+hSU5SMYkN0PGmGW6DfQpjmj1A8CA8uo3bshu9gTnVp7N/OTnNcXFIv
kWkuLUnfn+46TWhyJ+q0+sEMVxLM6+SPQ3Ie0g4UuxD32a/QW1WIxhKDJcPt7nEp
Wg+IQSlRiTkcoJXGRYth5FqY02z5+iHcocDjGszvXFqrhbNY7Dvok0Pglw4ON7E3
ftmPRaTLHiC4fKFK6yv6KDpcsBrbB3erGXsVJepjp+b4hKMOihXdLgeW1OChbnNA
3tPeyllbYUxc7BtsnkXNep4lDR5qNCVAPpMZsKpnAUtmLlFhrQmCm2J3fybfQmVt
qFBiMzQ49dEDE4Q0gQ0Z7DLJucc9e6zK7RDjBeF1J0/1JN8rrrbiavPhadWRSCZb
c+H1wGUK3jCBZLRKiOzjedDMG7p6hT5OWyztZ4nkdk6KpRkWVoa55rh+ulIGfg3w
MIA/aQJ8Za3G4RVPkwmRaI4eKovmYncHHqrpE8vwn/MY1Tnnu2T6Y8d5PX+TFOXK
uuJm7r6HmbMLaOGrDdd201507ISTSelli4PgKtS9fMm0BhfPQ29AtEtYKnhBT6Ub
WRIl3niDMLsEIjpHKeN/h6Z9w2d9vJXTB8Cweu85iHPXe8AeSf0HlZH/hpbLVQs7
3eD0Gp3ixzTxBRNOuquXIYWghL6NxHmigwpM3iyAF5zlQ9n6vvcU3yKqVsI5Pzby
pUXl3h69v9Exa0S1WvxAxCUOx0JaiqvMheQO+M+u86PRKt3k5Y2Rq1WHzUPtaDn1
Rzsdglx7l3qfd3Xkr0Oo53IE0LpeIGxT2NWr4avLXZQaQSIaeOpgq3NV/fx98g4u
LxC+HYyGxrOcc91gRwE4gJEeflgn5RRg0rJnk/Nda7mHzeVS+Jkh3waJsbEnnjmV
tRRTLOny74srshJ9/r4x2spmp9vJ1zfgoeNzRQMsx3QS2KR/dpVfQHccq33Em2yi
Ui7uOjiGlrXrsv4SVQYOqbzrj0bcqkJ1MImvy50mYzhA1bQQFqdW4ytIV0lA8CYS
X1Tb90KY1eH92u+QMj8LCsdesiM9cGzY9PsW80oomCfnrKgBVk7LW/pIdXWM8r5J
sawzD3RPQrz+DmnzG8vPRUll3lEMtNQRREoW1d1mb+n2BOUq7rcc5QKaDlGBM7VI
jWJH6vvHVayA4D3b8xS8Jvh0NH7olB3h9+ZbGBNLIQe/VNd1z4NiYz/3jZc0N0Vq
gC3B0CbUMwcXMN+VBYR/GWJFm7Pi6AZylCI2mTsDeLSuKO7rApLxhHQ03vBvZjdA
IrvO7MKw2CNuj++8SBHLKq4NTDYB+g3zMaBTonwPKqrbJErLhkho4dnKRlYzXpni
dlEjVj80XKd8sNOMOsktrqgzMX74R/Zwt+LpEkHpIswKHjNiEkbsxeYyN20H5nOk
nIuCZB+0YzEk7LjgpAl3k5Rhd0mpcFz3F/X9NiVV9tw98PD3dDh9to3EGz3MnIvC
ZzFdTy56aXFcPG9HortirFUu3hnTzBkaEIi8c5FZ8Ki2BFdvbNgnIML87UMNpA+U
1Ufg96SeMHXOZrMmhRmx0FW7NYjR0qbprRT00H1KsKEBRwqMv2mLLFDAvU/uX0Pr
Xr8EBduCWQPNU6v5DNCao+ALyD645cW7V17+RDmKkAIJk9GEWZH6R5MtaM+Arghw
jJLzRHRpR1NEYW83wZp07FPezbQTtOTPnbrunmQda89Y64BFJmCupiXZyDN1dOoM
pHXPsAJJBZbh78wg09oa6I1LOg1ns3DKEKkmTwY8y+bnrAaGhGXZXdBmPq6UhyOl
6Id9+djoxTW+Ll6XG0wg5Rke5RsIMvHmpmzdh9PTQwNNpcNcZqXi2ZBRC687PWhF
JE8yiKpFyAs1c3qaTsgwhYv0cXEmMvts7D0lXBhoqw/DXzQiIFMcVW6VqONA88Rh
IZurfMVpZQ2s6tEmzOQYziHP36IQYKoSgrzuK+JrER1XuIGVcDyk45ZU+86l1rMm
wXFogSGZlrhioP2htYaqK9aNTwa4586F4Ir/GBRKAMKceo9T+cuq9XleQjbaNv09
HpfwMmPktfXGViPTcR09bX8Bj1BUleDb2i12psdBuCymogfF4uj0EUqLyNH96Q+y
o4q36OxE4fvoAfLFKp2EIhWavVwnzEdlW31hNXreNAJnxJZjllfpHMnwB+cIf62Q
0C3+jv5gWDOcsrpMpVn8yFF7F2jmFj7aVKmhVH9tUX2fNlWBBEnLIovqAd9I+cXx
c7cEEYimAxZ3a+a27EJgRqtKefxv7FpQiIctJdHhp+UX2rJm7z6VaCMyxqK/ipPi
EuMY+zl8uXQRrw5HKvlzTF4us6q3vf007LlCnrK/wZzxaZcJ40eQU1gs+tV6KglC
0f+wFVubCWnpEvppZMHhAG1RLk3pBYj6+wPOBeNd1iFiKZs0FhP8Ev10AneQJFcI
x+7cZ5G0Od0D1GZwuqrFeyVSLSluwZci7qBbyD9V2wqNo2pq5bFjHW6+AbtW0+zJ
VyOTD/xzMKJTo+RH8DCyfk6Q88YAfr4IwRH00ZbnL7f/swo7Re4jzZLSb/dhH9u3
O7QU83XaRBFzZUX17c8AwQ0QKSf/VDTpMkPszQCsSOe2inlzBFx0r36pCojsGPqO
ATPqRxPPZGO71u+bhmtg7qTz1EKSY2J2nlibzFblxi1Of1RxeF04oozH9y++eFwH
aNMnc/Nz4edmvqBBzLNLCcRNJ6YhRwbF/ErjiYGkkzpYDZcYgMX/uD1Eve2CKI39
XGoWEPuzGblZOcGJQOQ2OiMMq0lyg9TEPRYuIsHtOKhkiNXvV6MWstDbIx0Vklkq
IqSREQALseJtKgvRdPILCuOUaui8o0S2X3DlKca3zd5z0BxiK/gR03LuWhN1cCaa
ATtClw0zSd4aKWuzxV8/AAy4IF/e6FbaBnK1jDOy0qo3m2UHQTpacii0OCZVMMdi
l358QYK7rrsX2kRS1zQ1NbvxVaKlEIX7lL60wpmnnfMFMc0zIYqt0ghuatc3I+5L
dr3p/BVyLd2PaNAOcF8TsuJ7pvAyqlzLTVSAQ86Lz9vy/luYJd3+lw6frAM/dHj7
wKmLsjduya8mE7txevVrIZUbhWgJXJ6rBy8iKCBu3havzgCc89vBTf53yIsHVP3/
WqV8KSW5fguJAR9f3g7CJss6umSS8o3yr9pmjqRVTIYtn2Ldx1hee5/KPuS9eedY
71cLNOCJaX1Ihrr1yFsTQ+ADOgT/o8opT7NJmybSHQ0cIg92tNvyCfYCCQFIhyNm
OCd06EWO31Lfx3HpKrXXPQHPQ6i2IQpLfRFCFa/YpX53yORs1+crbbzp+scPD4N4
tGUpRiLaABKnsHtdJru7PgIdazbegE2RXzk8RQFZbG/rmTbgnBfKiKVLLclaEe99
c0ZfoJRAnb0UiKNpRQFjhV8mqTeHU/raK3GlWTiyiDU56Ha35bG78CVvIxn08zDn
dn1q95HP2YywXIY8qu1E2LBbBhRz2U8/LfAVxA3C2He2SquQOVhV9eGZmUZkyuEh
Od3eFdAXV87XO/LqcQ1Utdh1GT++hDD9TbiRtUbbFSvzk6EiQ9lL17X98nFAbsct
M9kf3rnElKR3/aMMqdCPdjWtFzFgjGWRkvM0eR5FetdgSUKi4ZbN6wqq6hpIwWqF
Hy4WfLUFvp2N0/7QwNFtPlonFyXHDN8CoIXlj6ZbTMxv8TdE7juU+RslvjjbZ+So
TzCxcZwC2Qj6VGGQb5seeBZtYtj6L3ZE/eYEKRsE9OI+cHqMiuXa3fpQ+bwby4o1
2+SLpuG7NsJzfe/FGpV3qTfksn06tJng5pgb0O6KMH3LDeV17GxBfZ6NjgkUvto0
NQH8j9CNdXrIjDe1NHbBEkElYsDb3vL2zstlGs71/nHExG7HfKPospPzoHzhTHQA
f8USONz9lh9YpIVMBsrQVH376jyeSjfJ6cA8ahu0L4NT/HgB8tOJ7ZKime/rNSKH
ITw2baJyBBYYPiZUc5W/yYWZFrNLIyTe8wzwkyXwxal1Hld/irqdMAbHhZaLiPx4
xEuYnsOm+F4qNC7W9i35uKv/RxQs9YIagpL6yc7vR/F/LbyKSbPgrH7ElfzMIuFx
Or9lqJLAKIe6V7neBZVyIGssxKXSwsFZw2dBbRpJBmOVsPBM+Zoj4BLcD7myJNyy
kuE0H4JXeFNIqp8TZh4pJrJFH92zvmF61ehhKFgFVlZ8XYSYPWC1eJ8jNoS3WsKQ
xEbZT3YPMm8PT58k5fUSK7RwUFjcFo8npMR7FPcj7hFNMQ3nZAHpLTzkol3Jf3Cu
3lA3ZtLOMErUCPhe5sOb3RXwzxRxkDCzP9592jCHfoZp6tAAA6+z8DyEDQaIWYcC
TreYoxcVuTdzyDExLVCT/t82F4ii8IXLG46xh+mhDyDUVupSc/k92keST5kJInPh
0IovFrL3AcSkMk+7JA1OJrNa8Ksu6AsTRp59eqZpl8VHhYGPIkk+imHZeUHCP3K8
/+5SoqA33nGWqJLEkk/pHJJOU1axBxerS9xeXp1WMSA9IOxl8nUOziQjFkjI4OBg
uF/o6D2HI9UcWrxvGa5oAVhZTNIF/m0fm+IGFMPSDRxyxz1a45TK2ArBON420I7H
5it1cTRKFDJZpDbo6WuXEq5Oq4MZAlU+Jp79bnyoyIiSLalTWQlU70nePzj3MFzU
G2f6WwYRWQ0nuwVdVIviRWgZK3uRWbEk7eFGCwJSJOZ4WR2uXEwDC2hu+ee6rxkM
DvgvotbA/OF6jmVK5DBxYNqwySFbQDqxd1UJvSL8AkIeqjRB5aN0N8siGlYuDs/+
hRNT3RTW0P5C8nBeqSQ4h0h+HK8lsJrA73prhuLVLVc78lw4FvBMUdITAmL9XGhQ
E2Yjc+CyQOeCXjJJao208OJCRsRyTii3ZrVeeqne/Wst5lkULAXMEr4djfjIiq7E
QwIziBa6rAhmCZCTp/zpXqRSyXhjisOmZ9kY+CxVBc5S7zi2ZIsOlz/3gmCRLiMU
DYTsHistfuN3FQ4n+kM1EhN9WtpHh/AJ0TN2/iff3m2PIHEHpxdsmAFekF5lzBje
tVZaeTQkXHs+r/RJoMkw4I4mIU6I73iFFQbMEuIFQCJyiwZa+iAH0Jzl/649+JZE
QtvzKJgPkd4NFlwvgSglfC7WsCECwelwxEyFD2nCn1N9FWa3jceQOOg+26puV43k
ZDOk2UGX7yWnBtQgCzX8btNEvuL23ZKhwzMCOplxvlt7ggYoEoo+3gEMCCegxKoU
JuzcySjztSzWz7Fy5GqGZdW75nkLK9cZCWpzF/jh4VLxAELvTaC5nI594B/N1Qog
yb87BKxlDjizgkLO1o8c92CDlQ975amwjyYEmIL76DOBET52Rq3Is54vV4jiRqgO
a4o0H5+sMuJhUAC2XRGIYld/vO7EuV9hENt0aYCJ6V8B6BLqiDeyUtKlkIDKM2QT
jUeY3aLhWi4u4rRY7kd5X1d0iqmsnVADbV8Uw4qckdBeRQzPceY0ULnsR27QdqQ+
5IQpLXDFotRtJ5s0pI/7gYSpco6xWAr4igZmGuNO+xgPz/FkK3HUhtPxIm+XWO8B
0x6Cb87y5mSm5DDWUzHg0cUSZBx6uCfebOvgXtjMag+zI1e3Nx+cAQGrgxj0174J
zG1O5uw1CLFY8zW7LCrfp+FaoHGe1AFL37k5sgA2fa+CfLvPvaBABH9nplhVvdpL
g6qkMbeNp2LByoEpS1lClgN0pHWgLlcyyGbwt89ECaYXO37BnJ1EjgBMamK9R6kB
P44daFs5fJsa69m1CyFKTn1xJ2LcaoMlYTCWM9eT3N+T2iagjqIQaeOErLHqfBnQ
0yRJot4mTUydnWXj7eR+Vqfsr2bmbZEJBlV1F68wQBDAgndcqQP79UzY1gseA5yX
QzkLsReBXfmxENkbiGaoxpZq+0A6IZYtsRm4lZ+9BQ0RLgEQ1bSXGUr0I0++lnVs
GCkR6FyrQkSlCrlup093nzbGgL277CtuEK+gwuZFJH541weG8i80HPHzkAUaX0w8
otBSUDxYsGky6ryC9d7+R4tSlEBaKjP4lxrH51N9uclOmfMMAvF56QN1a651rXas
NGLsAYi8F/aCKoVo+BBwbDvb9uIIAHte9wPI+/dCG62bU5YpAzKhp45CzmP5Lj90
gTWlVhfwlVcO9Q0W0/mb9SpVRR1iJXtbHHaeFDecRPc6bkdboLo7GoB9ECf1JkbM
IC9s7cI0eQrwJ1Tv3u6xs47eRUIyuJz8R/0K8gUKuP8R+li5LfYCKm82rscJOzw5
mQufuNeJGrL5scSasSU24G5gF+MkD+m7Fxr39nuuOfwiURgclNUbN8HfJzXkTLjS
qL5XpfVjfjc9KPmXB39nN63XG0FoE4i+b3jIC3s/QlbjUWhF/hoT/E165wJK90/P
c8fTKDxRGPIDAn+wBCv+jhQsEeEA60w/ryHaNer8jnvFs9cFUzUaGQvCWglZiZXU
OSR/h/+9e61AV3xth0iqhUjCC76z9ECvsTSiPxBeAFoDM7XXV6jrdRjRnlQ1nTX2
cvaokuQj5ptlGKD9u1pEz02GzEU9M6y4i5iwOlniCuyxyhsmn7IO/x2E0j7C76Uo
yZx6+cTQNQIsNJvO8MeGcwXemqrjxNEjW6BQcTiEjwsPcBozdRUjOtycbNd6Ab/z
BJNzr/FVH3nJ9qp5zxN8GqlTwsacZNcLCFejcLI3IXjwRGVnCKFSdD55ie1OwK1k
TElA4pGU6SmF1tSMaZdPcXr5oiGlISdruChKZpK4t3hgpnKAQAMCkkoSsHgYQvYW
WkkAwR9lCXqBkBfT4aTcbqpkdl/YO8jT8R+663HvWs41YOfkVpzgb0poSV+KjxVG
0uuMfkHhJGeq1QlQYslKbUK7NI7tDB/YXu3d00Iqy82G+ns1WFuNFi52oHxnqRSl
ouKhzdjAHq1zrxNFMLAi7GWMaUxnm+o5wcJ83ZlLJG+MNLExLIAltLgGRe5aj4o8
1wwMASJf+I0pJBvBNYbQwDU1rKcVmBbnTJZm6fZpCAMWMjavnmcMFEJ6L0q1CQPv
96spKvZoYxmmpFawq6VrvQQxtmjEpupF3TXzkh+ioe0eSOmxg8n7EuAqBuRla6ls
x2Ep05qswwjSAMKWOgEhDQ/WQ3fyh73dsVxlS4BMH1sjFMEcYoCw0UzI/cyzf5xo
nN//sKDourkFpm3h/jY9mArgkQjT85b917Yy+o9D4XfqRqCzs316dqkdSgN0Z2U2
Wvda4P658mhGokgZoGxnSsMGGkeCqtxTqn55GltFsuXkstS5J7L64jOTFh7oMkug
d0Ip3HiAKfQHcEh16qU/wKz4868fpMdhP0347fwVbg7sykdQkZ9LPS3OrechGabL
+iGmtqf/hMtAEJEVnLcWV4b0fNglCOFzcXyj8xrrkahaALtDwKtLVCeuYjgWwAbw
xq1jC2cBvRAaHpfIW6jYYbFvrqXnNFF2gJNfh6Xo9mqVyKO9aAjKCZD7WqS/lqUd
nr8I4Z5alWOOAITmONzEBy70qk0hNFurji0m1G6+V6eQw2K2lEhsR14KkXim/B/+
wa111bvWliAb/NUWHvSHsqpxbRrLStETuejJbSWYiQ2YJD0Pf+7Apmi69OfgLlDe
9mwc2fZIKK7/DW2g6pqQqs7spxI/K/QUSeemOr6WlHIl8/QRPEYapj4HYi2Myz22
0JDvTiqqDMZeJxqmHX8DfSDocbljWtPEH8Uw3uQqUDEXs4XLwrpDZkmETFwq6p0p
DU0/Qoj2CnQaGsQG0IdS0Z3YFSZlr96gXrys5SmAUyaXiw/VZC2ZxXDY4th9mUDN
bTCQAal+27QNFvVJuzCrmRPrUbjtovLGojs5nfF5FF3uvhzEAz3rzWX7UDBl2VvU
qtpS7f/ndSf8hppuSz0GWdv53eg11+wnvsJzwSe766JkrPUgVjP9qUr23UJ62GbV
+z8SHPni68EA0TQnATeqnGGtNUaW/yUd0evwD6uosA8G+wDjR96d7jhxqeZ4t05h
SxxicBMv3Ovlh30Vn4fRV3aYw0KBv9DGR5f0qoD06G1OODnoqmyZ25WGKWoJbAph
5fR5KzuBKJDNXZMJua1HsewaH0P7w3uJM5bgnQALouC+MhWy3sjtVKvJ/5wDrWEy
POhdokXVGhQb/SNDbP6vbELtJMw/+SR2v2R6C/ZEGNfWcO2rIPBWONeSUVplk0Ud
dL7z+h2cV2q5HKjzflSvRx57NEKVaM7wbZXMCxefZRyjAtmVSVJZJbOKk6OVWRpE
xuwKJF1jV6bMVYwtW+GyBHAkci/NcR4f8g4sVKJggYP0Q/2cTve7VHIQ/rfuT58P
7yWZlZ+ovhxbHMkYgKsjigCmosvZQuKzN1dEAzV31on7k/Y1CfkzNN7Hg1mGN2Vb
RFJz33TRgXEF+As8HLD/BJeijktbWnaP/V8U9RHn0jl1mvhc48umggL58idKuZo8
edPUmfbYsogh5XfOBEvDUrFE5b0X+NgFX/ekzJsCFD5qFGjC8OA6wF1dxjMlCmME
T7ZUzX8/JUqoyIVZgCpFc8F1yUKDxULbPSBbBKTTzwOnQUfhV9EUgUkQ5UnwboGE
Bj715+QZ4kpjXN2bpWJz5m4yRhqZRRQ+1kqKu/wCqFSQu2LkeNlfkhQWFOr7OUTn
BVVlAJYNAG7Ht1zZMCbR8PPzp92WU1+JJpPMSRZfNxC+FwgRGzSqvPoCwoXBkSxN
JHr56hBfH+at5pwEH67hd8sj8felLNnpO+4AW3+lu1xHyiIcPUEMtYZ4VYCWoxzO
57tG2pvMj250q/1fq51nu6bB9AcpemLA+ThSM0IOvNBI1dyRI4j1hCJHq+rDYIVB
Q7waKSUyuPsqwOUfdrGvKP1ZAGpJet21iS/Mv5NxaPDAThtSDXNABpwsUA1/w0Be
0VswnIOxX4gYLpQ3/bXKUqX6YXBQuilO2E4xKz0tlJ9IMoM5bylfeQc0iQDF7tet
xfBDEQHmf7XhK3Ms110sNAvwMrAIUetQQmJoQDInCYk/Cgd6CMhbKVhd1ywINcxH
jM3y5TaZesn0TH+oOtznpdZMmPcD5+JPrIHT9DqziTeYbWNEWQCPPkMjB5RXiJHE
kYbMjeUlmFnpgheWPnW1QIWrEO3aoUd/RWfiTdWk/AOZYS8XCsqiMbvcwGGD96S3
5qRyJRHdxPBLvpyIKPSeRuSewZ+kFWLnJ1UvzzFm6ytOBQQp5PvCC+iHGg4fG+uH
2Emry+SNF7/WjKC6TEUKaILkNcZHFnh62BzBzxI8DlTeYcK1WqLstCGikqFfYW4I
Ze6xeEZkTwuGZOS7obSxrUQ/FBF45z1dfojHAPWZwKg4fYx+rZsto3jk8KWYc+VU
4a+21xZ8ZW5vIxdnJnWK1aMMGKDeoTkIuHSNq6DB/3WPq6q52MrNjJsLT/FATPaN
TXKadkXXhyc8pqTkgkKEC/ycwgtcd3KHmzXpfpu6qzhe8iiUZujSXURIRR26Zlhl
00RecO13f0AszYMigAESi6DyhUokM/aQj+35+8bTSVuvQYhP75brTnNzqEG/+cKj
ifJJT1tf3vt6poM/+bn2UQQHTeOhpTZYifkGaXsAXtipXTy+xG0Zrh/2pGoz2tG7
aTJwlEfXgZaFXYpu2y71cmCW8ctSNnllHgMmpBuc7ErAabr+89famkEC2p2QrIlk
oygeMnJ7rRJLUSOuOVNaV1hT73P4MxfPfXLN28PvbMECUr+3nJUSCARO2HKWSnuj
xCCpAKYqz65gi/G6aJWxRoTQFggH4BxDyAsDsoRBQiDvTWowZyAHgYg0jQOm5tQ2
YFsYfaYSTGATxuczK0XnGK1AzvUPdo5t2tq36pNvL7kUgNpkdSvdsDdZlK1L2zA+
w1styKy19QvpXdS2Uzu/teTwy9dOdOWtt70slJkqDIimcKEO1XGD/Z4vMzRfs/8b
ooMwMgYP9oP9pDm+mNqrfdYVf0/8JzJHCtHJIdgJlGXPJXowdhfEY6uSy9ejJgxZ
WFXM9l7hCPfHM8Vv9DO81C43R3MIkkmJyFuQOLoyCPpTaGu1I/qs1HtOSvCXjC0v
d+sBohJITv2PC6ildSrR0lafOvfhBYxS4IOm6Pty/ZBWWRUTtrJrDjL802Gat6FT
sX0Dy9pKFOx4mhzuQGThA/4gyJQ2Wt+XO4sjPeFnTNvJpzuePOP7gcNBlT/I+cKt
AJDfMzZSRV2kDlHQG+Us9WXgy9+LmbdKQuYGy2rtZT7xJ4DXYEs8gkHYaL6z46lz
OAIYtAh47tCXc8v270DoPmknM77NwJu8QtEOSpB+0i1f3zV8u+74KgX66rU5R62k
PIVgh8yKyV2WU9s9iXvV/Mu4jEZudYbB5jOVwOEOjzHo33mYfhkugXptmyVYXDDs
F02is0L5islkMib+1rpTYMCjHrMGz5EhdE8eoPCqiYLljsIoCencXWZMObAxX3t/
2fPu0xzNoBi+q8efcPQv86VW/CNerzIiS4MV7pyUGMRoDzcLycI+wp5PPD4/VdaZ
JRdb+gtMHUG/wHZneDs+u22PiaOYzrKrY2Iz+K7tllpmi9sK2W0dYUJDzEJsxR7I
IuaFnfSVsgQe2v5WZZpM27uPisyK4y9w0pp6MrK2k5uZH4Tl3bEtuPd/HP8OtS45
JhDppqLmNJpwZw8zNMvm02Uipv3lIMkW3mImILDyeb8w434WkUF8XHWpT3A6vIt2
CFR0D/PxEfPc7aXw0cO/oZFlI0LEb68knYl6qLzQ+tdMVZMLUWhYoRbyKocAOZSA
RIpD5a18hiPE5Ou5fyN3Gp/Do/rFDGyF73SKLOLO+TTSlJCSNXoeyczAmFmlWv+/
wmOBLX3jLVH93lA3npuiOx+vK/LChTTXUO7CRhuaXCwdl1KXUjjVI2hOh2nAS7/x
/XQX2YdC7MMcTnVGcC0nKyhdeNAeVO/SDyxRlKhctw6ar7nhgVNTL5wyOA4Lt3CE
npKimx8yVRX/Vwl68sb6y4WE5zdM+qXgSEKcZFCi4Ys3BPF+F8heHH95b+CPfhFf
ZPvrSkOfDePgKNm4fERE8TF7xZDHHzrUlEw+zEc3sjl2Cpe/9hQ3RlIMMgnr2YLn
J179+Te2A4+CpGbd9XYSWnqjBIU2pSyOv8x+Ue77imgCM/8zfsZqkvDPhgvVc7yo
O5x0sVd/kfCmDe2g7zy75hoXOHt9Jx+z/xdT7SFH/fgsBpEs8awVhNf0+FOE1/qY
sWazNh2jmWYSQ90UT47wmnTRmgXr+YY0xLoBzFPxWnD44QpI0B5FHSgQjZ789cD5
xnw4eCKo+BidCka3U/uPmTLtxUdmNGmIWBLT9E/dBN7Dt4ZO93Hpz8xAMcxhww2T
mwxdbieTAOKG+1q7D5CmmZxpjhWt1vK2JMhk6hl4pjdAXdXhoGG4fcF6mD3mJqhh
NAcrG7RXTASEAtR02Xab2+uYcVWr7jdAzCv0SOOA78Rjb5iUAEfG4bd+joSHpuid
KEqWFs/0I1os4ndDIke+KPof2NQyW1BdeSYXHPRKtrlVjDPpPyOEWkYoxLQQXw/I
JmOlSXgJY8EBc2F+k9j1Z1muMLFn42+2mJLNgDmVFvc/44Tsym5Z29IAP1Ug2xYX
g8rlDG/5f1wr4RUc+OaoJaDfWifya2K1SA17pqNLzRWyZONZtSm41q7jAo9/33Ir
czm/1be3VMBo0hEqeip8veZ0Xog0OqDHOciRkcW6kvPmdhK4tkDCclf4SEIQS+01
GAby+ROoASaXYnmvIDkMhhBGfMiJStg5Ux4fR6ZEHGa1VkmqVUIgIAXp9/PyxH9j
aU12L+dB9G9fpg1oqprEJsX7Zqoa46ywGjtgpCUDiP4CVMsQJMbMxahpgZxpL7//
xWSm9gI2H9LQs2+3J+f/MgED/KGQbBG73qY012UqjPw74Ch6kamTy1tM0FtWUwbt
VzOBG721EgNGqJXZU+IbWhSatINZWT+DAJpoBiWUK4HiMkjrjLpOQwmSfxMsk8nX
tL6AQ7K9f+dLKFsWYxLMXxDCKqi4lWKRDflYeOQavxzWtGxpKWstAlUziEgs5riT
bwmz7iEfY19+xYIQ+ELmHUdedrAceCRlX3Q76NH7W8SuNb1zB4WsG5lWj6K2BPSk
JnfJLlUwTIAC9rJZnYndarlljihEABuPuGWnpp1btEcnK1WqShNc1JJF9Xif1ZeX
1SN5TQyU5E2ItXvRFjgQrgipOjptHaqsCeVLu9T+cU+5Du5ifBlZcGOVhEfhvEzn
tpAQnW9OhdPk+FV4ddrw3kIATFh5ur4E+8RYuZetw42OKIAdUqn7sdn9AGSpVxvK
3jk7JVgol4khIlWm5wuYXG+rcDjiYNDhI5HaZ+OTzaADkOcd5puHtH9/rdGfaSK2
AuqikCMZOXqFWHJlCoaFJ5t9gVUlYG21S3P7aUE8sTFDXif9CZAr6BftteYkvkxa
G2h2E4Lz98F0QDNZ1sCGYtrQ3jcncComtKHSpsNHLemNjA2aEzLnGTDSBBQcZkew
z+5OqJxvubIAnGSW8IuxAxRH/2iJ8oOsam7lBjinVlR1uMGpLQ93INMa3MNkrkOG
CRpAliUEQjK+s5DC3wc5txSQfFHT5U4fVbOtexLFhIWxN/CUAdv/ARnpBEhE+eHn
eax+kUzqWteml9gqn7MWixUcgAqk31RH8O8SD4LrQblTP1KTBtGSAiUMvZqGkEM6
M3Fbitkl6SynJN1G/kkp4DFrIpYQ1u49cqkQLWVRmwyjpaXkvU27XPXrpoqhtNbX
y4prHUU6eRUBJpqPMyAI0SBWioP0gsXMQLzGWwIHS3oJ1rinucfyeiA9r1KvlHIP
S3DVIZmZCuM4IFSHYD0h0Z9LQ0yq03l0kJUwric0Oxwokk85Z29JuDZLoShM/T4K
M+RMkTnyUPH/Ubq9okuovIByUKaJbRycBSDZ+yiX53OUqkfPZhWNaDsWyJDlU970
wfd28vWtPfhoBGFsNTKlOjg296hTMK7NhTw+jgAG6530QrvQBs1zlkOXri0bsv8S
RTUP9URb0Y2VMDLcPAdNlySAkGEs+lvioVjDmgvhIs+a/cV0KAIhCyRgUI17dq7S
h8J0pjuo5RHnkGrQx6Yis242iFR68QIXx98cYZ6Pu3MgrhRLFQkeiejOwkzboxz6
r1J4MFuGBS7qAmw+vqVDTAD6ZEcSp16Cxq8Qgr6n4oQeRkM7lpp/h60Yoo+8v306
SbzidH6FE6jJ2PkJNGmp8x7deHYrcPzl11svO+PvmclyL6h+PPhRancJ84M9bNMP
X7Oe073TQ6oUeVgaYqtDoqvD8JdIWKWvvrahvIt/og8=
`pragma protect end_protected
