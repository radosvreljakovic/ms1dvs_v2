// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AAtM4sRCefhMxgTOPbSABR++4r06FWSPfzsI3H+gpbyMbZmOoWbm6KKA8wbYBW0X
9Ng7olZGDFobmzWpkjLC1N90yRxov9gbT/tMvdQJCxsN09aQVrOW1R349Y1RGFeH
080ltZiNPeMJxeT1UZfAiu1DU0V6V1ZQV6aglx7DK4M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17648)
9GuiaMaIINnyCO3wbMGzPaNpi+lTpbtfZUaHrVfMBFm0SsV7iL2DlZ/i5BqLEqt0
MbLSlCAXyRhp6msRKIC6Le+pI5wBWaqrNahZxBBGsPmN/do7El1aR42JDFcI7K7X
icMaXu1lS7rLd+Q7rChZmFAZk5N+2I8oLE/62VjQPHWq6yJj74ARBgrJdK4Ntc1/
uHanHDHzzPV8d7p6lzNtavlJdy6R1/mAHxJmTdjvhYPY962m8RHYan0gixc26rUE
HxEHcgdikzw9tc9vJAFMi1rzDUtmN1L+Mocddiv1AyCmj/BcntHOcNC3VoAU4bz7
K1JQU8UOfPGC6ABW+zdQajhL8whFtn9RjGT3j7La6xnxUEqv4bT/OUKTNmCUVU5r
7QaApzC5ti0Qz+P48CLWU9wCT/9YwOSKTgILIF45jGXihe1kAz0OGBCshJtt5JPR
LKPaByu8kFN+AJAJDlnlfPM5M0A0aLjy4yDlknkO7in0too08+EGgXF9sKCrLON8
yVclTO59bH5AY7iRGJOtEMSROp5oyUrEohnFdZerGNlxgVGcKXBBDbg12c5M/EOu
Pt5tNH02ydydWALxTNaSPN24Ayf6O3oe1j+eKTokDxhpVGPOSOdDjiAhIhc4uYCY
CaweNLz0CFOiRfwbDUNVtk1mrkdEjzX6Qv9mPD4kZkIjEfW+utwrXrXQ4HAkGeTb
zDMm5QPvWB5O5opSRf2lIYuvQFJWa+plUb+ns3SjXB93zNsBA1NZvMJ8BYKaPtSC
uxVVKEpmYH2ILHoD3HwViMym1pE7tSvqhg6MRFPRCc00XU4nYwnvGWxQyWsB1f0/
ujVo29FM+8UIf+QarR7yGsUhFjWMP9uy6JRwGz/puFRvl58v6/K0zUcj5zixtRFJ
kbS4JE3uY3LNvYpFiF2EuzTY0vVsqgsGTwHMsri+mjPBOKzcxyVtbDAteBMflv/C
a1youXuGKJzQqbfrlGnL2U5HxRkzXEvnmjHui0iwm/gDONk8eBOD/WXe/cYwRfM6
7BCFbq5krGMgZECpaajRZKp5rNouPuj4/NHXM8Tf6GowNBkrlEIv+SAk3epKZw9G
czX3irOWdxVCqx9alBeBFQMd0P6mZnXLjkWm+QSUVQmO6r/ZAJIc58rK20oeCv4d
ZBKlmba/5s3Ul2uWGISW8keyGJPaoA2sO1CN8iW5Np1JyZmxNlZEVB+eTw4QG5mX
L4BYHq8PIcb+g5GaW0p0/cDs71lclVNnyyhAnbwAmWjCNsPmrfIQk/pggVNxDSsx
HwgyqbEjqjRsYBiqKeIkVAEYAw7oXvLMdmBi9OvNwOVWSFNJcfLbYfxht7IlFSqC
CNRRKk/hRESHLcwcuhAQh9MBf01BBZTegOf+3q+oKb7oV4rlCeSt9safL+lwtT9G
x+T+IzxT1AxPbInoJLkouoMCnuuzmte9ft7BYcY5k23ABZJ0ztW0laoiMF6AKyxB
rS0+8hC9OanmdYZMiUg22lqSRA72U2rt8//tFdIgktUag30bBwlcXlFEIZZBnv1r
lgbs0QU2r8Pqc87blNBi0/e/fkzpSFHPfMxUlmPUmFLQ/QLQNPo4wcyZQuKc2X3w
RuW3vEWoPKVf9GFcKW2Pc25fVJRA1mfQpH0aJJ6hPlAec41sks6dckkOUxOG4X+2
8qF0bK+EBIrK3mJlVAh5WFB7M6gQNodIoANmlBKV5ubLprWTTDaC5NbIFOm7F5kz
QzGKN5VAQtNlGvddgwW/prnhoPWxo8tO5x8ue7mwPxoHz4CLDN7jy3VH2nYw4Kpy
oCA1mcfj/kGKZ5Fjwco2Ys03PbivG/0VsRTFuiz9Qgvaa7RUUT1FUnwgAwaZ/KCW
pgfKgi1nSohaxBuNwM1HKr2Kw9knV1Om3YA7uigtpXzCZgu6fG1PnV3X3qKuLHqN
zneGv0uzb/uUw0KXMhVASrA+XsfEOZoiVCwYo3cT2ZMDaiVN8ovoUcRaBgQmXUh3
Rt35IaA+rMcFugkfQZL/AC0PaBctA8CVJNQwBMiyiaaA+JzUU3w+xsmlN295Cuqh
qIOpzlhd4+87yS3RWZ0m2NIrg8xsy8CpDpYBopCGPRJkIUOZe96pWHu2d1e5HDlL
4oSvgm2S47quqhAKIPoQxwg+7/Fm6n5HuNz1vxDZRfUsRx0ndthWJ/nhPtml04RS
SxUPAHdUtVCiZSGiUYcvw8cRV4fl+lAsJVtbbNfrYKMR9eA4s5sNLll4hDI03pSw
MMdmC2TAnY11jlWqcRjjbSFMsqZbyfBUNMfyxpBAE+UxHwhXpmdRaI+sVq/D/ngv
ONlnxw9QTobrSUZtRAwc5pOy6VW5ChxveRTZA7JvXJUGoTf2HfxZitsPaYihDGGD
e/e51uUyMG6qWq1pbM2dj9pWIjQv6YUDrn891vxhIWGOP90v+i9hbTOm0rqVC3d/
ng1s889vxTJzmhHKd1aK+GPQsYYEq2lSLTsyQvBK7h8fWeAbDIKm55PtcIwAf8al
qj8WMFCjdQLgNg7aXjqJZoaBjz6g9eMq7UE4B5iSNoK8K40n28q2hJwYkLmOw5Gd
vhNJxyUUYt/PvTrINVJaXvy48+AoOEwDuvKEfVL5+U+nWAjYa5L7dS/34lhAitQW
zGYfAS08wNdZmWn/TEr1K7G6hQwLwLOaKzaKa9fY5LYpjkWk9qFJuwuSL6G70tUO
wZFlKRrrtzGsNYYRB0b/8aDxgU5zC/R4tZALnKEvtEKVDGJRXLAB2XJh0Cpu1/Wn
h+I5lC+SJeWzxcMCKdRpJglXbN3a9IAo37xMvXMOvQqvZXcPq6u6o9MyAmI16xo1
+2FaGgsfqOKQWc7B4kbBGxbewkHQ4DJYQ15UxhcURKhLUZvzoRuWw4vmiyrEpIyA
ocMuoKRFGNSg1f5RcT/CmuHE7h2zO36xJdAgijZkxkZ3nbJaYe+K5YoLmB5Wg1FY
3u4Fc/S1Ce/Thtie1oU0YT4bGP1FgOWjMUQ+RfH7J5Xd+g+k4B7DTkspHv5rVm3o
bptFr5Lgtv/LPu95U2SrvPZkZDCH2SfOJew8pXi5xOaWCEGKvcI9542B3Q0sVmZc
RrMiPTUqLjSAk+uoivarZVwAVoQVk4bu1I/Ii1sOIUEgrXDgGdkwk91mhOWmoMWF
EeK+URDGTcg9u+sFuJDOuyIdJxG18uYvGdy6eCld0GoiypUFSDorU/6O9BOYj1kQ
zUEq49M9Lb0mFMAtxWaF1gbhXEvyFe5wm0vqgd/9N+LrdCkGHaOT8Nv2Va0dViNG
p0wwFpXVKscsKFNSROIBbp+kfmXkLePI85We/BOrF+KpiTCmXmrEEW5/MqxS16KZ
pk/J6YrWz7AaQtk/tHFh1bgrpFO9SLN1g5Ott+D4jESLirqTydK/Uw8Vh3wvQIBV
IxK6Tz0YCEtKt8DETTK8A+9ppnIaPAIBFz33E4e4FULezf+Lp9CmQGkDywjyOjN3
KIFWxZMv/rr3YZisHiz/Ldq283+QToqqSncUCPZ7hztNPssf+ogZx2UtXzzFwO8y
BsenQqkVKxp/DFEb9sjJ4Y9cflafnTTWI04WpWAdoNB3JHgzuSs6S3tlY7DEl6eA
l9t0tZBmpusifv3pwUasLTDxz82CiHRYTWE4uHQRzclRebhtxtmlrBr7O2zgLn3l
Q6efkN+h2VWuGjLaMzHr9GQMtzmmkmx2vmdSMk0AnTt7QMVU96PR+h2NXfcpvXhC
btdA/Q12l2YuK0IOVQm/C6wiWCyPtLvvi3mmCAcRsu4OM3FgJZTOybyW9lg3l/xP
aosthVr4I+u7oucjNn1cr8vzBGhom9OcdzS9l1+D+YS+mEUac+/SR9kyPggEOz+W
qh2MHAkAF7gTVKVYSm/3oDC9yMvpzDwe9iiU/UIPc53SmYp3dNvxVXcOfwk8AXOj
bUiOt+rGvTZjf5EyQpJ5tEwtkfzuy22h38pVzpO4eyTIB27LNIejE6LteAOFXZub
BGCi3ICaGOHrRBa/FxImplPa1x0wYDlbGZhLNNkBACR/GiheGf3zzZ51P5cHjhrP
WGSLymUXGYSh1A+uYfgKCNo3tok0nPZRdal5+ftnjxnTbcalBeOAhwtN872StIQh
1vGLh5OtMr6Y1IN0Zx9xs07MAWxjDzAyhGk3Dxy9guSQXvHoT12ZJ0Itbcnc+XYc
MUTo1NZmI3uN9N/FIeSUStLcEWheJ1BDYAAOclSunFO7a72lFnoE7Us1tPdeERz8
GChpg++NTAeOCp9wkkK4F7NZnmOQjWksVxrFCKJcuqLFfTF00Wb0T60QKemp0UzE
8yScfsCFJGzZv5PLKlVRmhce72t+9LmsSXHkWuLv4iBMvQWdlv/z4H1bx9t0xfAS
1fgzyS8Fhzl2cNdvjYctx89NP8OoZzUAawUSwT44T5glgx0NTGfjvHYww7cePYkr
wjTaQ81p1H4HYloqriRO9cZ3LUeUTa3ifbe+hAu7Yc5V0C81jIGYIapwu8rd3S1H
UFf0HRPKcd82JKTPm3Uh0KfV+QJ+uXsIOiSfZv9DKDuYipCQqQL/hvOpXTnJBmqq
hx/h4zkr6KNQmM8gT+FEyRzS/cVjcng1q0hDrH0FlczMMagMEsz180bshV7plt4F
x0d68b3wiRUDRsqIHsvZfsE1Hj2+ixim76W9nvjLAci2Nwl+HPpo9Tc//YrlPEVD
OS+fLBe/zfA61hYw2I1S+hOmWQ4fz2wEMM3KLyj13zXUZ3wmU0wmnca1KFBbLD0M
g1HkaNk7JXYt8U5cnRfY+tL6HuYCx9ULEKrKZ81Zh82thdF9NcnKZEx2yqAA7L+3
lB4lyC2M6zFxhkclG5OobnrceSu3owNfvwpuF3XDv1rSvu0bQyz3Fe1nGWG8RFsu
5USaekX6R8GmHTXVmFcSEBTmbGZHBKMg0lVVY0HUBAt2xUkVNmQq/98ZXttGZfaI
3c1beBDxpIUGnh2GDfKbV01C/mPqI6e3cjuptR0mamrvF5mX3k3j5l1YjOGY2KQF
ByKkVDyhAJqsMJqbYrlHeJlzV5DSlDdtBkS+hTRgyy4h0Dfb4TjlKyZM3zNQHQ2d
7wkI9klDkCV/8gphdI49ap2EXYCp88zDdCofoCYR8Vl3AzsBKUJtTWkDxU5T7RQh
TVNC5aAkofHULvs3huhc5eturI9xkmpt/7/iCeLdevztmL388sBe2KgJZ0CbQpwa
na8tOoT7S+GWy0Ff1s+99x36/Jc4KQk/ebVsJDLHruN6n/lvpY4IOWJU6Qc35Sgx
DQwAU6GkDD8QFRBYKkPDwVOVuPOW0AsdkuqV4ferKcZooKA8pM/C6J2S702d2ZZk
QdqQQodN+8b6v783LrQlz/zttU+pZ7zmatNjDfinKQcpY9CF2iRFkP5WTukWgQCT
aT6zbGpQZu8Uq6+x4yX6Pq8iK140wpD6m6ioPI8TOf8sSu4aL7K+igkaulRCJ85Y
a3WL+9TgLNTr6v35wqca6+Qs+zEWm7c07qLDfR9GVsRvZjxdp1sDYJLugclYmCej
qRtU/UxQXYwsX5jwwUYUdMvPBJddREMAPRHnLJcOMYbKEbffZJLTf5v7/akPuVgY
rq/uO0msxKaBX+Z+EdHr+LRV8nROXAiYh6DlRDNyqTgbp9yK19uiAnd5KnEj/Xc7
r+bi0dbsMa3HShofv18MOpYC8UeQjjMgN54vHsZ5uHXYSrZ3fep9YOlmazyGUHWs
WWQcrtM8m3YOQzRImUMQ1zClnF2ItMJAge1jb+7WTPxHOf8xMQ3OZNSCaaE89W7+
qq84UP9rxpOeAXHA0jl9RkJb+tUcW4668uSSLlm19mDVl+hsaocaqmzaPJWWKG5e
EbZOieZEfAPv3Y0GeVfziO/g3c4tKeX8QKMoGhfrBOL/XxsMS2j/Qyka8ItumObj
e4/T31PKsclj48VkE4W1LGq6G0MkS2qoHRtjPFUX0F3s3XXSdhRnW5CVV7xr4UuA
Z9PgAEtKde5y5agaa0FwuwDEFFVYcTYrMfYGSReYl4cuvBDD+Kpe/CxKQoPVChTI
eAGERXdfQdf9/+FKxWFdsQwIK+Tvzu20rj3E1tbuoiB3kGnEaO2kbkrapU0aHChk
GnNuuSYd5fni+/uzcNqBd+21/4wppqOCEaTuYMOaqysX5/jK4gJLpBkK7+Vp2Dbb
aeQxjdFQrqAx7yyNyGyfmKSr9JcBb17d+ihSau1SQJF4qfU1FFBhr2I4H0tVP0lc
AY3YWQ65bDsMLOOXpZPktP/A2miHa/PUixrRa3z+HaL0AXbda+MHeo1J5uM9ITdA
Jg36/Oj+BnEe56EpSalviu3QUUBgxnrS9Q8BmuCowKFSEWUYuin/C8M4Av/z4No0
efd8s4MDw6GAojiK21h71t6C7uIrtEdmF5XgBoohvHAvSe6mCqibW6ImwZv37r/9
jOBoE3y5dAh7e6OueFmzrek/zFNa602/LcVnjAbhz3vqPzw6Go0fPiy7FVBhNoex
C7tEIYLI6jWQ179UAbemrL8zdDoV+Y8rIzzUPkj+TGV75zwTqiykLwDyNw5Cld8W
ppJTtZov/cCLi6h+iMv5i4NYWF2gp1RDF48o2jcQB61YpuingyupldNgEks8fZLC
70Jaom2LhvoDf1L44bS7yVSInkA/9G3S1gNCQjTCHMPIuKy0bNJdSDYAYnxedxnG
1Qbp+v8NfKl+DduaZViDH1a02dmtMiL8V6PvriKB8abH6cmNWokc5qjZkjZEBiYJ
YtwVeHzMvk8XD/5dJxu6Iv9WLjvs/UF2O7oaNyqUWFPCmxCSrotS/LWDfPNUA6ou
mQ26zflOlQZF9cu94IJ51zAcoH6bP87rEK1Il7XTJJ0paY4vV+wWDXmBHnVHuBOA
zyDYJAgFhFqwXURAAcF6aOERrTq0/UMjLZanXFu7fGqP3iU7f/7i/6fdHb8cBQwU
Mugg/A/mIUfj6CaBdXCR9qEwMOSckZ8LV0rZb4cgh9++Xc7FPL8oYeaQmbXUk5wU
pI36F5AB0yUGG/RkMezpCZLni9rWxIEe02KoJNK0PGu6piRphHJInjnNmIaK+RuQ
6kMsnDEYjXCFzbtsyZ9DDLkPQPgP1xo9+sU3bmSbMO73Uoj6+VCY0yTi7mYuifwI
L1C9zplAHVVrsiXDJuFD1BesgFxVgLnDZbWCDtca18vmAsE1LaRC3QRwLMRX0a6l
cP3Qy2CBiSnOIvBHLkjHnuCrUvQueOHFHTyaYSG1Kzh9mIb+GoLdWseWisKIw7Fc
Hv626VSpWkeCXWR/gCyaSBy2vXDmQ5d5FAcRLJ1pWluafKIzTh3e/lEyJPwgziL7
zi85LHkrGL1RVKeKnH0F0bmiHnmbnVodafCXMK1iiIvqC1mNkdeHCka1HyeQG+kh
EaLZ1sm1NU4OhQuJ4ZrH+nKLODbByux3hdqOgH5+nWpdpVOvJA8j8ZuzVBNAIs33
3H+83IKf/MmC/0yE9xDEPGLh/3Tvw4R4pgAlphOf26bYC4HzyvUfieCZhzTbL9e4
X98E9fYHAHO7Z1twB/MtL35QTrHVphEveQaybzXMqzZoh6xQs8S45msXtdLDfwn0
ncq38FfcfqecIQcD3mv9ktxgOfegEKqz+cJ6xouLS/zOncQvCTta8uj6aDokXNqa
CGWTy5lBvxqBW0fb8MfkTo1lV6CZh5C4Oe3Mo7rXJ0Mj5817TTSnPe2tVMjVB+J7
a+pYV7VHujal4kC/XcSBqpl6xbkPR9MOeTz6X3RlnjZALEcGYzzT1oKgm0Z8mt/6
H/IIvup8Z8jDDKBinVJxjxzma8H4lNW0mymInQBtFBL4oZELgVCKWTeVPNrkMuNl
y2KP3gNHXlyqwrSLBlXVt3ISMXLrZoRGba6KmHUvTjABfuSCzHyml9UXTEhU0sHr
/xkMRHvwz+K2kl73vg+fqOL6HCrA612G6h51AIby4OvU3U0F1ZuD9MKC/WcIljNx
hVD+SXT6Z6DN0hhEUFXbFbuBdq3KWPSeCfLPZ/7Dcp7QkmgDAG/SVXxsjw1uTg1s
MVoFJMo4Gw5fF0vw+aMOBUfnUpWuWJa8yAXdH4YiWZqfD5HKFwITmw3nE/lNElc7
dOo3NzsbkIPjXjNv2cvxTMBF5y32dctbdQ3QEdjWUC7x33824/hZ4/Arp2Jf7D/j
Aw8E7ItlhQYBrxwS2fOJJaGcJmsFFmNnx0wsL8HdmW4X4cCjcpCFHwClMIvn0C8P
C/J5Oc/Xr8Xrn3Edf7bjcewgMJWvL4WXvnLCAV5nJmTuGozouXr3FbynPsV7jkY0
DfBf7n4HYQLj6nDrCEmi0dviKGiqFNM4UQ5QtXio+nWVyBjH7yRTUBUQL/0b4GkL
NVrpR285+RF8UG69Br0odiO1NqWLb1pAf08umgIWqg+eYHMSKGX4s3ZKvq8bI1yj
EmD/awZj9yI1ZC3qS8Vfsh2H9YvCJqzGRsK8V7BPg4UFjsV7FYrg2xK2YAiYZ06n
rZso3h9bwmaNoxVlNISxFo0pYg8Sne9rLOYgPJ5taw7uvjzcm8NF4HztykQUTmBG
FzxgGon+msKhBe+eL9BK7Px8I5VIfT+Wt+i1gyv69jFl2WNqjWV8CrJ/iNh1pt1A
bHHar1pAXdLK+VKov2nxzBRhSHAo3sNlXZduW2DsX8v3DwxUJ/b7pfsLJadBbh2u
4kBe8zTxDtVf7Y1A5SE0sWUWAjS/xsjT83NrxRAqMKDGQNJsgViRJFeNYmt+9Jub
7g54/e4TN1t8tmHlNRUUT8URFslPtWo2rjKCFb3UzptyAxvRZqFrsTEM39U6i8z+
c3WAqUOSj/7f86tiIqfuLtSvFXvlQd4trq6MgyihE3Tq5JcSY4ygKdLTjN6G9/Y/
SHNDbto1xIPaLYsPA2h5X2OROjdvh13B1wEQM0s/w6dS7M3a1G1wEWPWsSpkHY0U
K93JU9FcrhggP5JLuF9UpCAxjiq297ssXjBaQ2lieoEQWpgvFJ6nIejvx5YgQ97J
NbxNPouIXmNXsqtj3H+KGuT21/FIiw0daPgJAvYfyXCsPxoVguIdNT53fPyAfDVt
YBB8iG2fYFt4ZJMTTGgxVgD+RmK6fAEMcyMqqaazWbodGwrVuuGvqVK1HaDGLugI
9d4ONdkl42ltJOyflIJ0gJRGzEpX01IwHWfe62qOFd30jPR5Axuj74ypMn8825+T
VIG3gOllfJ4NlYufgO6Ksy+Tz8quh/vz3hOuEZgI8olFIBZmMDbydmtffeSVjUwm
8E59r1UZb3pD0G17bGqyox9ueUVwPj/BuHTGHGfG4LWR3TVyUS9hMkELo+sE2JAn
fD1iQdWlob/Oo50ItRxFzCGphQdi0Tp0vySDE7P4Ltq+i2ZZcL9AkeTBKFy30IiY
RyUo72bnyBo2NJ0CV+WjVIgum8Kg4z/RjbTyjEUExCE2tcqgiywiUgEie+TBItyy
D5737fGwMo0MIHe9xnp7Hq92nWKbWvlQ7oVRuPOekm9OVkkx+CUynUPjCMoRP4yU
9lPvGblGrNKzAk1q5OOdZxa0hgyWFzWlf0o6kVHYLSsj9KfbLNBAeV2VnBgSisDP
X0BE51Z2+n9TKfYta91jgSsOKS4KFSfiBQvHcN618fut4NcmmBkTYJekE2m/8BYt
AZkGAgJ8q7siz/PLFa/m6ym9G7+R1FO0XaMB9ncqzklyyIGLofmYGxRu3HdqCnGS
6QfkLoeLgt/q80kTDXuYUviDY0RnL/nnXBuF1VwmUg0JTg9J/9muZ81rKREviRA0
yDZqKonzj6MqAl3QDA/xpcmJ0+SR6UUF4l8Ic6ils5FUDF9yzTuUxM0GArYbHxpp
fzXaVeb3CUA1pN+vlJKzC2ElNwFrBQzkFWWweNL3cnbnCoN+PPpls+o/LNkpTx/j
shuiHQ+cMr9c64N3Cpkg/OeJjpnz4dlXHPIjAP7WGQWhBVpOqrcySwuEgJr43mH2
NT3STaT/zUtpAncMhg/U6FolmHBBbwef+sahA6KufQLvQn1ora6RjzSBvX62lA6B
tuT5evZXtFwIFxG36XkgdpVWXKOdnrYExUhFoRGiNDBkfRKhmcgeGbd3VLwhWZOt
NgZhlCyNxwMt4uyB40hfp8Fp/0SI/zKIumhpf49we86cMc+Ol4Ch6UoMgreRp2gO
2kGZPeCxnU18C/uq6gog/wp/ogZI8eVjMOaMu4lP/weMNi6LGmM1HvzMcX81mN1c
sxseIY7vKXUbWdUM/km2XHN/RV0ONAoborN1RHSIGV/7oSMZ68ARDDup/hr7GeIv
fil8oVBBY3d8X0apjmHzFrAw0jfj1b7QllK69i0npXE4le5f0IkYTFjyWlKalJQV
U3AgvE/An6vnKHmrI/BzjmwyGXQJlOcWjirsG7nQjUNcjan9xcJrriZy1r1yvxCh
fGbMde6VTO2ZikzsbX2u4Rd/GS7nrrIyjS2PJ9Ht5Kra1dW4quCc3Xz/OxDthArW
n+2UJuXKeqO4eSS7DZodaddWsTSnygeZAy9+nRWNDbfdO2o2DjelrMBJeNJxes3X
fBwgy8HVrp52MLgyL+Kj6hfa7NNT8WYKOJeLg+M3pba8hIfpbUPxWajXjIeFTFye
fvSDiqMuQoOej+eeJgnTwfbAFofkvVeCXnTsIcafuKedjPx50Dph7hUrNDvrpIOS
1/F/diWNp7XIux/lBI+1c5wMWxlBzrAzbCBGODyN+yzRa9t5PZJ3kBcXwcX/OK7W
cw1MjeX6KvNUqLIgGq9iaIZfcQTOpzLOL8FiMK5yx6eXVl7mmnaRAvhMn7sndJvr
Go/R/eHaDBsS72kuaFwx05apDVuq7lZ8Z8YhOqBvBFNfUfO4P+uswRKNwerTsRqv
Ki2HAHBnuherkiPbC6QsNu3ZSjKp7ODaD9q9gRLoBpz8g2Qkxe8CA6/Z9rNKcnCy
xNuzv5Hv0RJZ6qgp9LIVmXHIFyRC2TVyRLrJAFSW3amyOMSrPnJA2BZqKDvHKzr0
WqX+Cw+yhHOz6bQ9KAK3dRP9L5CTXHNBa3BhSOpR9RgUm2QX8OJY9zXHm9MqnXM+
II0IUifj3XQiMWtad1AuR/FZmJ5AfE92K02hMrg1C61JAzGMMGxOwGp6Dwntc1tu
FK5PbMlakZ4YoCti/61fUJD1znJf1Y+GYGfVwXRvP2tEvmiHh1gNAr3piPYaCbVp
SESI1tCN9dO9u7Esi4kyE/126V+xGXzFsoQ8+lG+06JEpexQBMgdCNL63TEM869b
zrvXQqZObz4DwONaXqfHAxStTmk23c//rjMg/a5IZLehhu3fzl2Jg/qfrIbVGH3f
beJN8CjmJEUD6DM80NkXCh602MeeHu8tyOQATZugUj9fi7DN9grx1JdoLZ/kTW94
m9Y+zYAz+6vWCBgXq6EyNjI4bJ689UMPo7LBCN0FUNQbFgw7KSHcTQAgvdddoNUD
K72InkFpgmYFdiVc2e8N6LclpTtEpnZs0Zz8Q76DAJo9024uUMtnePoXo8YIR26z
fGV/luM1KBbZRV88j12cA8cm7eIwEDpMn7ZYI/6MNSw6Y2rM4wI2M55/Aq/L3QLP
WLdNhFRMha9jJR3AK1ML0kEtQwvKI/SYO2M1epgwVcCmtffYv4NX78j3utkqjL0s
rGp3KdIUBIwb78jmK45cPBW80gRZP/qgP0wqM4pmnbUhfxNcafzqo7BM3wySyExe
A2gVH45rY2cFH/bdrTiwhn1kmKfdmhkaFN2o9o+6X8TchVRzQpgrWuuYBQsS7mo4
IQIqwudFwodctwPTBiz+XVa6UpG+MVUcdFBM93iMSuENrKq5GvaHM11np1bgupsH
QWD4O6lZ7OQ6hjRZEE4EiPj5pUHJXLoLF4bGT1Bh2BkY3oo50vv/aGlsPUQ7aW24
WlCxer2Xuu2L+8Nm0XLCPWBfsCpPPLFR/YQcLZavX9EGz355B79sQv1DScqPyMxC
3LYTJfAtme8j3hXNmdOWDVQGLhpcSsoD+7HEWeMkIRPysHM6zyN0+uVSwtXacarY
xjQtziMi5ajqoNA4HXo9Q/KoSPbi4DUsL4EAUHIPR5MCAh7tdGU3yyJUth1/Sk7d
0xRAPlTa7dsiNNOF4AfpN4pCM0Z/EAAo4UEbL4IvoChULNQn/gk8bpJNge/XazmD
dB+u2fmgN70zq1UKxIZDbeirTZuMtd1cGUkDpjjzEsNxgLe4xRuU9YS5VXJAQRkl
E1ibVpAFpblOYfLWcbfCgtedj1fOCEWRj0T1qXFuKAbieMR2o+QFw1HxAJr+JXKC
iEClxrBTwmGNr/rlUoSoDI+H/lCxo3l9JLX5sq08HWANsQFnF5JUL2MyvL02m4OH
HTGO1djU9QRAdp40XO8oeLdi4nhDQZcyqb5d21mdDdGFXiTfSlga60mvLNsexRxi
efKn3q8fTC3/iC8fP0e55UUGYY1CPiOohcCr1RhTGbihdZwsMFhmuawh0fA4iDHX
KjBfoD5xxLQZ/3kig0G3lkdgYrOgj8WvfdtRtIJakwkEGwlbYcA0+pCWS6ltQY83
VurXNbzIzcfS97VVL8o/lL/P3G2pmNTPOXTPwSO5BRACmP5g2XEPD1mbD+6CFBHa
0jEq9dDsYjDcCpJwf1z9xwsnM0D+YegE3aZL5Xx60pbkF5ujk/t6U+21quNZAoGq
omrD6HvJDTC7n9slHjzWUiflfM3s5Do+e42hWZYdsro02DMgleDuVzKZ/Oo/fP1r
gPtj7rjZolxHDfJY3AlHQmHsx3a6Jz9SfXv+kPepBI0Zh+WMWyUGfV68kAyNaJsO
WWTGwk3W7GlooiIJCc56082FxX5L0ejtIyfqUfp0/G5yVQXFSFny/W3s0pYfBvC5
/ZGhUlbwifkypeKxpGr0q1ZzWEFtZHjv5/lidUfX4qN/175GmjlZPYguByI9SE6T
8dHuxpkwV5dFxfMJUjmjH54Zqk02YzAusGgrbOMOvRJgjknmEaM+ZAxuwu+MwyA3
1brPWDLEvfW/1aApy0nQB+hWRwgLtR0zgDFE1U0DSrpKvf1SG0XG4g67K88aRzD1
AKia5iCi3AvNNPUYlfyZZH9gTKUI13xvbJgZ+gZnUQaDWosuup6jujcqfijQE4Dc
bxB7rRW79q7ztwWWmLtrCNAy03pYEd79k/q1kY0E514ZgYkxto+OQ98KOYxfKJeK
pZpUQqHzmg7hlT4wJYNFTZPS1QemXkxod+ujxCmZcdMj8z+w4zaSeLM7qnbs8eaS
m5DQKRSL2Qrb6wISLkvzJJc+Ouo/QMgda+Nx9JvwaG2zSWH31vSfXGAyigGl2WDf
bCpMhG17Fx6SkYG0YItmM2acTx8uhr1v0ROi+G+RQ3XHcQZQbl1BNlMDtys99m1P
Kt9P66wRHPYR8Zo45fSAEodvlXaQ4w5B7KFYsjIfsiCySe9wmbiwKUvYsivjl51E
4Hq8A19ypy5oHcGC41Lrm6pYsPZwOBssrYCcPivquLbEaMmdLZFaeYRSK0JzYszm
FsejbRoqDEVUkvyPAJZFmNQQmT/AipT9YI+dwtlTUuZjGmKrWrsviawXqpuhUWl4
pZZkqwlyu5X8Q4D5PIDPntC/CqghjqajbQaxT+kCTPwh23YIwXpFMNvOCCLZkE8z
y41+rMP7pm2am7Pns5Q2fWmrFyIqUH6HzwN4yzoeYM97PliifB35ynejJ6ORNlHo
lo2v0uqBFI58eSQTRdNNlUIw/V3F+Rz88TflvL+o+VQPHLRdBWpd1OMVQeoUzU+v
x3M1HoEs5IW/cGxBIgR2xW69maC5zVB32JwwWpRZM1ypWMSGIVmZPzPA1BVc8zx6
1QzDCV3ZoZJBzgH6Ju/Db6JzsiY/4YF+eKbNCU3ZPsmE9AMm/dJiOp/RjdXbHG0/
Y5WkxXyI/T5X5bsARmAK8Sn5QQHuE17mEYsi9+PYZYeBSXPLTmWH7SmNvabDtas5
thhS2WmWIm4Luh9teJvToh1kQs0joIxkTOt4PfZ/HDh3TBNpftUY0TLURcvgZzPR
zLAId1ByCIKVKpbw/ArLaDUMJvpjQ/QaDVjbbdQR+hXkf5OdOOszqkMoGuN/a+yg
fG5oDTyabE+YsM822HFbM4veU2NTsrDdGneBlJ9p32RPdKxnSCNOsHzFGA7gTq5/
IG05ScNn3jQo3XLK/yiWvum+PbH0eizTwTtrLG+WYSIw3EKmtSodlba2bMr4cp2J
A9ku+JtrlHJ+C/1W1Hx6zVKGS9pdPUafncNsFzMUIfNzq+oTdf6Bzl79RCie5YMu
S4EfdSEj2Ekd6Gm319m9y5zPRdNFw+poO7oFY4YE0UqjZf+DdfPVhhOTTfC1Ta7f
JV743HNjNem+xl/JB1ftlJ7NYn4+UD54TuizIPzUQE1/wWhmJ91WWh8XogZvp1Kt
v6VIpV63ivqoIng848zDewLBh4rIU+KliBKaDSWCh9LHWZeTWVgdscULKoHe6R/G
nFnck/wR50eTwvB3zdpgf9Vd/pI+dykEo15CysGr/KnsCezLgAxi1nM7l2qs/Wx5
Kvsonrtk2GCAxueG2xUa/wWTWcjU1c8M5SAqgGTlUhOkp/cbE74Ry8FmqVmm3O0e
9ENAUkC/xife86L94rimKO+tcJzlEK2Wqe6ySxioTKfNO4lDFxX5RspMqyI5YJ/G
Vfhyhh1+JvU3iI+i6+8ODm3eLcmuHfBZJVfwdNzeofppWnTg048Hv/YOCl8C4nbt
FghoCA7lIM3Kjjis6XR6/dPUBlrHlHy8yXqnNovOlpRNbVNBhb0GIa20ibX7HxVJ
rc2ZsIe1007ocSlkczaEaXt57c1sYP2FnCPtAl204Poh+xdzHAfUaqFDVed4u0EY
xSV2CRpOX9w0ulpwiRrB6/uI9mmGNhSEvbQbRMd79qJl0naIa9gET9cu1Ob6suX+
deFOew8neWWlqF+JPBSpNpSTHCSqkj/EGCutXA+WqHkgnLwaJ3TAUKW/dXQvuCUQ
ZsG03tPVachMwjaeWjjNHSCFFpAM97etlx2DnaG2qgjRLTQoENzhCU2IyOhRzw/1
uIweRWiJOCixxVDQU/k6VJnp5ixIAZDhPSewXUoYsVRgNb/AYS+P+TqxQWeVe0iT
qK6KDzo2I3wYGyPnYpLXTzn2gsQemq1FEN9OeIj7JJjha1JnfYinjI1nmvDciQK6
Ud3wtdY9e7nIvOlr/pkkdZC1gEjPk60uJCuC6Ysb8+FLZcljYUdnw9wDbLCUYFZI
a6HUziMEFlRNUQEyRM5z1HlCW6aY+RBArb/xYIPe4lacCuxDjqyOWqxgc6ExKhqI
DRB3Jea5O2KywsERRxwGT7yBHKWTczYi9Ye0OCxk7ThbjRtGmsRABO4yhX8Au9Hc
ryKMR3EfpxscfOXYG+OT0RrgwOqMHB0zGymwqCxpoIlGwQUTpEViSsarddddpHfe
0u9s8FYoL0OIowthB5prHUmHA4godNSfizUIIebIo8Ou/derHk8ZVzYXn1gOrn/6
BSJ5KwO6sJ9ZbQuswcyrAXK29tNge04QAkyrKGOuKxRiVEcfDzreRYY635OpT9+A
wYkSV2+gxTwJo7cWEqCwW8b4A5WXIGLkR9tnhVbhEC9AVw/lFhoD7+R8bS34VFa9
X4QWsCYw5v/QcfvQtOPH0eaYlVTT1atusf64/Edw0SV2jKu0Y01/BhjwRgJXgLQK
c3mKMIhusAT/FsJvrTV4TD6jFzLCPK5utoutdDA3y7I4BzlAwgdZd/J2UJCG7rST
gsE4CVSivlN956tdWaDCE1LMrWG5t6OiuzHvbn6T9u25uo40/mUIU6T0AZ9LL5gw
X6wmDxIhsSJxGrQ/ntaHwjV3K8EeWyxpc0yAXZbaPbmM4f4N6zvfjrLdrfS6l1Wx
Ee3212EZwtTiQYwxPR5ybw6tMxjWAtKh8MPMWXveHUNyAhFu0/cqicrFJukrWpnJ
BS6pdH9VpXUFrWpT8vxmlclDdgvzW27tWrnv8bnT2coM1sroM9BcHWGDaSnIxDnG
5VPO1GnT8LMgHU++mea7Bt7TMgwBVmXxLpO/N3OTpiwks2kWQBCy5lMQQkTxYN4i
nUDtxcVAU+aBZYpis02L7YXC/v1PzAgFCLgV+NlTOmGBTebMHcqSsoTBVDFNTr9N
eduCONecudWic0mWVTSgtGxG6gfby5qa6UHBGi3SfU5w5C4Y2qyTklhp30nIUWQP
CeRzMg+7aZRGQjTU5sNWoPvDMNtc+RILDj0DQuhbVPOXZxH6vgeM1gEL7l+3trKd
Oie1jkbQbYfaeyWORbpq4aB9el3Y8fuPydSjmIwxSJYM6ooWD7ERgZV3ZmhPbHiK
ymeNyA3uqb7IvTueYYv0AakJqiJB4jsDHXDRsIKF/N6LiruHFExI6zTczGN2eXoM
39jJv796aIurgNwiE1zO0T9Uub2DYa3Q+RfxJ7v5Dv+l2WewsSwoOPPXprBoon1V
JF/3pZuH+yeElAnFn2a7maIpZ2xAn0L0zF0rdMHyw1P/uW+6x9fOSRWZUfHenHZI
5D2i5imO8+qkw0MpcpJCGqncmcU6grbY/9T47yGrlOoABAg41VQDyKRl/9ofFOzx
F3Ol6rflXPJVP1mIHNXEZnibqn5f9kv7eugBNYo9MWTzMa7lTAAAHupgCgRl6YrV
Kg8MeDjk69eD0ygq+/GkY+aIdn1CceBE20pdv+/AeP5I/sieAMCkngRmuSE/k7Ic
MSaeGogNfXB7j8KcmVVa4dBuoy4+uNoVo+u8SaIR5vjduUV85zIiGZYTF7YhU2v5
ymADWwLTB0W8Ave7vDNkwWIRLJ/cbF5o/9LAEGYijuc7OxxSKD5/+tkH0XWPUmZI
LxHt8lx5TRiUTNYV1naoimJa2IYHiPIN5QzoVNdmxlbFENnag+kJcnoDXqcKOdgd
ln9oZBWolhrcK+c/LGbDpjGDK1iuOaZ5M51TFj7VVyYOxyXo8hpsXpKaskwIygA2
hAgyxp9iG27QOvOk0jabNfTBFkemNtAtY8Yg2BGuDroVshMssAdzLitKlIu22f07
/s+4dv970LlfxAcOc5uYBE/LQMFxvWOthXkF4p4QeVln3mnfEJIeYu37z6SYK/0L
8r58q4fq9WfIu03nYlKHGi5+nyxqvb/MTl25l3M1rI3Ou6utWI0srXwu1Ff7luoo
0fQ7BOiGtjNNMbyI3TspJ985CgtKPUUrjYPrykIAJJr6datmiuUGp8u50nAGUO0M
hrmo5GJgF/ntCugKuU6Ne0KSLxLC+si6XUh6GHdQl7YfIBUM48oZOXYYd3CGdgsA
hSrVoO9lYpz/nlWL02Wig17v52JbbLQWUNyAW/JxcIvBGuWecEggSEsMdgqrxcLB
XDSudVstiEgBHYmOL7BSr21vUHzO8C04uife9M94lc1HwKT5mnXgBGhsnmlTfOxK
vp9RUvEiAR6hpHqGsr9i0V4IduDT+c6pILZf1TA7DGq+AH/kFqHd2uw40lTKoFcN
uI6FW4PH759uge9yB63pmh9LA9sJIXiUjuqwELFVFvu2jfeWQEe9uNkhKaXNiNEj
3VtZONx2VsKoWEaLyFXV6dLKVW0tggtc+xNdUa4ZyNs3doqMBnyjIQXm8AdV4G0d
7QvKnEHPrJTmMPT/HH7Hy2jxeSSNLQ4xQ+hITsKG5lT7ra9EzcHT6UGOQeuk/kbI
cIZq0oIqwOgTzK1jcVL5daJbwWrKSuiPdDOywLEeZyaQ+vmoyLi0ZGlLZudh1IGh
pIviI0h+txAY9DOazb2eNHpgYOdI+mSOqq6vlU1Gqctk+1Ph2fYDgo3ZApqa+MEo
rDy020pD6rsFszdpnGd3z4Fm78WFauhpI7kf10tmOBHvpZPI3ivsILzWEwniJetS
ab1qdV3D7FVNf8TajJ1Udp/8+Pq2fCiepCqs8XFhXnUdZyLNUuG5dQJNdcIm1DpO
Dtx0JWuRHZm1caGxpmuYhYz6ZjFIIJlfxP+Fn+IGNBDFY/vncHiB1OYFE7Gt2HVw
Gc8rjt1+tCaigeOc6NPTlfp+dWpNKMlpvuO2PWRPuGzGM5cgZgU2Y/JMu+ZjF5QT
Trx46j6JUETDT7k8NcEae4nT6fV2tufUB0Ifr6aghdt5j0OUwpHyphwPRlFwxgvn
i5HnCSUwudunc2FRoMkqCjNl9IxiwbBcarcS9+/UlEwT+v1wVY0QYfPSEqQp4K6t
Db7/iCgI8FbvxN24+bRyMEvaB9Tuvo4KdphTU2irsiWAiRoW+TDHOO1vWlhI69fP
MUYwx3iyVrPH458Yuvb9HThpJoYakJIQCeJV/2ggXR6ntdqum/YOeD4YFqprvWJo
fdaFSOvzMTQV4p1Xf41EfZeNrXItHDZ2OrpSfne+1N/GoxkM63L3B1AcsFFrgt6m
Gsj+1521Eu/TeECaZoKdDpZD1vcHLIiyyEns821WziFzVuBufNcqvSFB0QVHLPzO
T0J7GqGDuGYbQwuZ8gCCfkYm7gbQSZgJTFIvogtghgKST9Jfoeb7cDqBVTFQgyPt
uhSZKW8U9HRiA1k+nNibxsiAJNAWLZWayhU09qTcUO72oYJbDqTaLgBGrcpaQ+KR
/313BUJdQdPjCt1gJAls7ZEhoz0H9kBH+xEVKJXZOpxdGbQeyBVRk65M+5uvEA65
R61lIAIv1uhfjsBAVWqaI7gd7skW/8cICHzkW0DRPdud+I8jOSrjmzAEA5J85Mkp
gGA+bTLtpwx9W/Lpfy8rPK33uFWNa5skQ5MoHG9ILKcpwkawT4PBoRoh88IgAFYb
LsnzMhQhVEonGeuiiGij0Ggq0ve8FeqYyBd3eFUgMlxUf7D47AoBddaPWq4oP1dB
S6WelM0XFvypLDi5rd442tRgL4XGWBpDH8QURwx3KjcOtNo1lEFnLzco7i/uy/iB
RifQ3jw93inOV1buNzFdC4xYDr3zvYADkUScOFN0+Et31m9EFKyPhweJZZcI2OSN
LLL4HADVvrfCUcGes8xF/IOH+MHqYrppOI9+4F6w0ESIX0ubtq/zPXrZTH5HR9qs
f5UJi/M+wDP+W3WH5ZUs9eTx9i3W80luFov5PR2EQ1SsPL33jSFwBNScnHomFqXb
wvqYM32Wc23KL8Y6R1E6NXFJRAQ1GEgUwjodPPU9KoFqSEa3B8ZFnblf7Mv/9DFd
pQ2/8PKA9rFpEi8CkNW5QeNcyOqvSLLISbHCwclQ7qBWNwg4u1JZRwntbzadBU/i
wTl66qmwE5+rg08qGymC3Fx87l8P9IsyiBSJlJO4DkQYQXOf0EJsju1qdlpRUiLd
vAkhwXAmE7aAWmmoFu7E0qqyWCzHkypE+KRdVFEws+T4RCkCKXxqIp2S/lWxq5IN
/tTM9J4RNwTEc9p0QkpJJPqrNlWPCTav0MYH7kAP34r3f9QLk8ezNle6wFqUDoOv
NqUwSR+RbfyIgtJ/9EkxIfogBG/Ze4NjeC0dv+984xHSZR1wmSuvyoWmRu9mHE7I
kWyXxmAnKb0Fyft6uOgQt5+YsnB0OwRr7AOjf8zi5MOgFgO6CwCqQmRo7agfZfKY
t0LltmVrs+dqvlMlVKi9BkA6J6Rym4R84AWIhu0CpqhJDCI1gQTnmyItuidzqkTO
bKHuLaGxHpbPECQ4xvnna48haHMz4OEvJeokKJbfCY/gLrAQR3pSJmfGYE7xZYun
aBBPGcdH5rH7+jye3cpxYA4h2wpF05aBLMA+tLhNH355NQhMtXnSj87J5rU81pAL
YodnhJDUqirNEzJT9zNZcFeVfH8zkGKSSQvgBcQ0y+DSQIYe1eT5VKnaKBIEcoya
Dwg247inHS8xsIq8HDQy8lggs5ySO5kMl17R3PcnOCYL5kZmhZvXIyBOLobfRTJw
zymx1fNPaljStzsnCVNoJJvmIbmEOSxvbJfN/tPaaEuBsKdyYf23F/MzSkhnNx0q
N6fiUyIzRjWEG5iY8F+NUTnd1fkCjHvvNbJJaX3HBtR78Jgb2IDQv1bfeuqoVfEe
S9pF+85VaHVHD/l2FAEbGefghcNgMnP8VB5n95cszCj1My2qIlQNBKaRl09xS8PR
Z3703rttCdQlpq7ch+5E1+/fWIo0/IQVyQp0E1rihJ3n6mZ2rP2LsJ16ipoM0DHf
lN0hB86P57x3Gipl9E0WFq608TmPpQg5pYXPsl14Lq3S0Mik7YaQ55OCgU/a5oQv
dONf4NugWjx8N3AdvzBfspzo/aINF6OvYnTIulYv4HhHKaRkeTKcVqK8My9tSPzY
VPpga3AGH3iPG5WRerME4a6PvV7Oc5d9fzT4Inn0P6/pdChc7FQPTI3SZhNupggu
TF1kGVsR9KLtx49lY0yoHzD7k3F3TpessEDN1GZoSI9+unAzoTQsBuWtj8N7n7Zx
n2fW63qA48P9DCD4ucZSutGC5I2+5S60eoo6Dzd3JaZkUAAeeks/bqJ3HPwZj4FJ
/c7PUFp6Uo/aZwi2j9SOlxux1Rba/Qi5Kdda6s42xiI3oLetLvFOsiQZoyoTRCSx
mhHnr7ToF0GX82t1i3qiZRqklxyGib/sUOt4WCUsaCs8hnrTlR9UNFfLQ9OjkI2I
hYPGd3dr7s+zj9dzHF5FkVOKf/pkVKCVJCOJL/DUJJx1AWQb/JhBMR/FR6kTD3Ag
p4cFJaLxvDTYXDYS+1sztl/Xdpy5Kf5CtQwBTfvGgOFf51b8A/UZRA16Hk9uxjP1
yH51jJ0E8KSb+v05lYP7iIKwIoC4kTjnWM6tRB9w/zKd68En5ZRrU1pHrTiMW/qo
giEuVbiOxvQHJEuJLp1LbQLWKP2M852Rdf4Zp52TAUT0i6F0giUwZjeQzcw+Ih+h
Fm5cbSlN7lrkhaFmyGRQ/U9VQzuo/ybncGwr2en5DWmocqRFETT7fGa/zPmD69DX
KseHqsrbdzgMiiU20tgrBXbzXIiz7Czhdq7/y5SJOw5TE4MXKYv2vkaXl2GQiRab
we3w7kgH8OTiTDWyGexbrazX51cmc9ZoxyGLDj93SIq+d5+5MhoDnJDov5vSzRjn
ez5xvsAtPU3E/7CdNNZZZ/aTDHnsvOu1ry9o/MKFgOEokc8NR6dDMK3+NAliEJXZ
Fcf371fPI1wMXjVqMQdl+T00WUB2n8bjO1h2OmOKHvpbd5ujzAubA/x0aiEK/jWm
NtFk711Q9G+ftjNIkve3JSS6Qb9Ap2ZZJ4jm7omE1fUNthMqhJP3YpTuU7jFDRd5
koRjoTIYZVJ3UJE08o9OoVg5XDcKCW4P3mBiB3W3F51jFUtOujHNI+Si1Lv6BNCh
oDqpSsGpO6fjB5mnx2CX+CjCRY7ao9AbmraBWrD3wnpzT/RWPxrwxtOuiz6wiMdB
p8ctTFYvAHecefpH9skmOyQlGWEX6za5QQvybz84LSwLVlCLUxB0BSay7j+hA+3S
RByFnCH0K2jiBEQF2brEZFxa8XQAE3Jn29yt5XLATazzn9nPxkQH5j6a7LoHLoGl
SZGh7EwY00xNNf0JWhDzQlf0BObOh6p3F/n5ApJojpdd2Bsslv5Nfhvr9YuZhAIS
x870VA5elbiI6ctx7SMuhArb/KJB2V97qmw4hAplNXE9/0ih9nuBYwIbPIzZwLDh
8XrLfVeWKPgF/Rq102Sn9zslGaowLqekKbdleooLzut2c9Y4ix7NTSRTdngzXhgl
oFRvfxrotYfeEuqxfT7ISJWMyWA0hXV78F8H0tKu66yl0QpUMl1aAPEMI2N+JL4O
A8z3w6KDlfaq+7birdDQezj/TdclC6HtpOHZEVz0ehFUvMyVQidVpJPPGeR/VK1g
x5cxu7NBgh4dmR9BahxeBJA7Uzt8qJPDyK+t6r3/8j+pOBKz9Srlb6Fdhy6e8zfe
6LdNb30hfeDtbWKToydh9AxhIMD2kIc614hmFix2pC0s2P/BGNWc0O8DcurWzCtU
fI5DfgQaqmB6g9PrPDw4o+k06+l3siLHi+qSObAe+4T+xsTUh/AJrVQaCvD5DfQr
jcIPJeMsW4YhSW1lakUa8HbY2kyE18Y8Nz8rQABIuwDeWjtQhYiNqhS652lSynsj
UiDGRLSm5n79Dm4r4ZzSL/YknjhniDf6LYLAv10rHNPE42YjkjatPNWGlh0Sg6bC
kyNRKgzzA7n38jayWPxWiDUjqt9bGm6QCAGZJbgAVxYb/xFt8YZqntSwoaXMh4LE
Girf4nKeiEM0LywyoOaLrTaNZCbOeLW2mYDorb+iy8dL4+BrpaL5DXA9F5xeM5g6
4STAp6FDFlnFdJggAVBNL1dnJnsAGOMy1UlLKNywlFQPNhOOYif4+o4pVjFe4c5f
ao4mSCiB8cSPwhxkf3Q0AOys+UrWKnWAAXWFRFaQInMlns6E9KpFYe2EWFRxn+68
zQlE7hXPSKaWKjRZ905jb5ufkELTs9xom7aQec5yl8oNxb147RLj5nvf3t82hs/O
C/Uth9Me040cf70mSIC4nrfre5iWeCMuXFDIvmNgqNP3ykFUqTKjCl7rRa1EHMp5
3BPVqwuStxtXyN8y/r66rI5St/ugrxn7USq20hGO/ZueJMELhlsrAvLBSmi80iKg
ED0TuwNZKJ9cfMrOX5ynm21xO4WhMCMJZV3M/3TMmmpY45CFAwbK4DhT8OO1FONw
UbDj+1SZhDni1tnm98B0KjLP6/wrkUfh9xvlTi9FOxnfeEG+gpGxo1aSXAzGTEL9
a0OIA+0Umg3nJCo0eY1FtM8bs4gG3L1/l/eQbf0/o4p58jVT4B+PjTudpLzoGiV7
712vwLluN0R854Mq4Pu4gh9ry4z4+Gd2wi0M9j89+NPgD+Z7HLBzTbBOLlRX4dT/
6xBhrJM1TiRkD2S5NlxiXXnmrVpCcF7PVkbezuL2y9h05kOQ1HwNPMnsT1F2tFTd
5SNZ9qx/2wWrsO8uaut1RW9KPPkn+PZlbM7MmqAjlXkFVCIRfkCUBpjGpkePaSgR
VdZ8mXhtUnx1T+tI9+5vMviJk7VOl93eU66/JkoQEFNZJzM53o4dLJXkzjd5O6nV
yfoVDZ4h27RHAohVUBrprwgBgKt1HmDye+PEkECOTBb9BM/KH37XACVLLtSLvR5b
r0RflSkUd9cACtIIByrUUGXsB/g2nHLFZcyigViGFOvxklbe0VLXzJVop5fKHH4c
74G5wyRwnUK9mlQyc+n8nsIzF7KJ12rDr7YJcOzSkUim5NFAynvgLBxCk4spphpq
xFoYKMHySz5sYVWE0GPzgh1dSloSHFO2rG9dX8AuIfBywa1UpfELuwZcnJJjYNTT
hMNzyWEuY8kgiOqvbMmtuvJ/1LlB4f50HtsyZ+97dwFPfdbWq9vdS5GuOYa2jL05
1WR6f8Yka7DDWebwADdXup95p6K2CnHTGO1cLVejAbT83K/kYfTdy39nnCWuRiXc
zGXBjO0w1aUyNyFeolmwAktTW73zQgdw+FyOEfSyVUGmQ398/hgmfEGetLLG0VLb
so7YgFNJj3r7a4krPUpQGtNOnQrDYrn0XKWJ/XdFIpqoTojsEi595fC0Lsmo6zVf
gspMz8wXGeCgdr6ZDaB0G8iWZn8iW0+bTYK0fet0aGhvb1Qp2oQM+tGpRB5Rc5eu
slxqmcwz2TUmF/ijTeilKvSrosWpWFX9q1Wmfnh1PYI=
`pragma protect end_protected
