// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tUWj+uPpubiSz26tfIalYcur/IxWIXJoLCpIRjnJ7ybey/ERbAzphx2rMBbdAZJ6uC7oG8u6YcuO
/guY2E5ZH6NhNN+PDoElQ1E/0EpnViOMKyUvVX5qwlWpPvbexITyjjsG+8WiN9ldD5krGtnTavRC
zzIwhR5KEW0HpH0Rh0G72vvfP34yi8tyQ11HQSPA2eG+yI/Jzdee/adUEdGW3AqGolOBMsxdFXYp
Pd579S9cb/HqQzxADbElKiPTtNcC39Mjbi7kO21pkdg62DUESNKPZ84+PzW7fkAfcQJ0cq9U1SJZ
0/Mc+sEpGJWWdKZw2BcB2RBwXUvjEBlo7EYT9w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hhTugFkjK+pv2mdVEpUOPHfpatHHHw+LBXV4NuhUvPqnSGSn2D5eeaYOTEsGl/LwXki2lSCxK/YZ
jBibraCu4B1b91DUkd6kOfEgfATWbb+PHg7CeY7xaZ6uHKMTq2JwqaGbladhiDoO9faR4PFhzmJE
7FvA76pesmD3ZiZQG3mCId4T1uLUAaAGObFgSkF6t1Bmj6ubxn6sPxs+C6g3rVpKQiqDx5D0V97u
kA6zqyLjKrq98CMrv9UBUrlDhyVDhWfPSGwruf6U1VIY+Me5nin+csuDgqwFCm6UIxXNW0E/ZTYE
i5i+dWro3dR3L289ncgSZLqVitkznqawxUXUi8xXXFR4XmJYSFJgD2rTyDPwv17EyYbopQ4y2dgK
U21aM9/b9IQ5Kzv5RvDVoB7li56brTlEhqoTB8OLCBzReTx4LKK5LjFn1aTwQ8CJ/wkApnYPT4vh
CLFDzbC6nWPIKVhHBgm+TLPlnLpM0jX4NkG0T8nDbIxGIwpEccxs4I1ZRqQsgTz/TuAOH5ivfLeE
c9Sudx7nmQ75/gBESkrMNQRZDzZ2oC+3yyW/8lqb858dZvkRfU+o9tJ5nkEFQiVpdwSZvsXycgPQ
KC2381MeQw4v6IftWKUdhg3vLXZI9Mf57J644DYfLsqR6/fNVURJe7IFerE3K+7IMi61hBZEAGY6
djWUMyQ3lnJm476QoXUl51bRCs8O0U4mdCCZ+DO8VleHrW6jWI4Xx5G9GgdijY1v00X+ywG471c8
IpRGMOawAlmjTgWU3HlawEcA9kT8WI39bFRBa4GROG05K/YacXJ1ecS/36BEKoYmFWz3bKbC7Te3
d6ofyG0YOTdOawkhetsxdp7pW/S3RF6YxCyTda+VOBWHA5LdO9Dxjomr65F3CdkdUY856KQptSjE
hJsgGr4nMJjWYjjvmFUCwJ5fBWW5mJfiyYrr4oKAu/c7V0QxwT+ygdwGtWhUBNOrn3kBklMyBC2m
0rZ83EgcRHPeJm+KZTOvcC7VrdO6iYQIa0U5JNAGO1WzggrbBPU0pWOkptFZS3kRYRNozCM0q2mK
xLd3ZdZhANCoAkM+6GJC4GDJ3JpwS36qsWf8/KFBVj6mQUzvG1eoymF6UJ6W7tOYtwcJZdTF2iWB
4q7/0f7ZDyW4iRFyu5E1kG6r0fIScq2kzfnLqGIe4TY0d+6xLLMJZ08NA5zcPN4jgKM4Zm5Ya0rq
f2Ko/glecQI74hq0LBslPH1XwF16kw/TY/vMcZtKwE63gT09qBbe+2d1qdTTf1IYN5JjFIl8SZpk
CveRy3n9GgD4OR9UDqrc4m0UKB5HvrHKQdzPLjb8ZRGa6AtjuRrfdAJNx7BLjgr7cliyc1lfLZqm
aZwTPfwHFUdLII7cCm2avHSLClwAFFoZO70k1pDhLPOPss0j3rA+hpfx+ASyv33CcZMet/1QRkrw
E0tQD8kpTMJ+1mfdlxOCjMRdshFiagDAIO1L+PGziNnaNdHh0wU2bGokO8gXOkTobXjVUgcVzzI+
cURf+sULj37s/DDPCEU495DOdHgmNTvvaIBZPkH+L3EYepkaKv3QToXraNqe5iB8pZDm/EIIHxrK
IeNH/CuqcZIjrKT+RV71VaQyjlqcYkrbSRJtROEiB3TauA3kJwGY0rK0QLcYDo2Tim1HWO092rkV
IrF6iwZ9mpItUDnNfnav/vca/Qfqlzmr7PjaSu4FOq+C4GTbc9bmtVZ5hdSw6hKY0KqudhOsJ2Bc
yAzdlXeEIzejZpsbmGAOIfdIG7R9U8w+ZC00BsYblMHLLOK2cjsJAwUHNt4qtEAB/cr0APfflCuw
uCOkBgoD2bA0C+qH5ge3LeuUnC8TmJUWiO9SvGL1ZxkziZuUCSmuq+v8/X4TgvfxGIuk5GZadc+E
H8CIDSOA7PngXWGOn0ZDB7qkPkHEWLPlKrJ3GOrU6ZZOm619wOR8AjSwssQzNiVAXtwdtTp5ANsV
VhhKRDVGHMjrX0ZvQNwbK9Mz3yOXicm8ywXc9IHgIvAo66339M520X5SPu3sIYJGf7mTeRmDq6Ja
pHjiex2mnZCWpw12p4p/5eBM4A6KvN6Qp3l7at97j7YNl9mHsAk0LS658uCAlA9N3N1kzdeR39sa
3ops+YYZgiAtjLfEHTsM7HkkMgAuOhgiR/odzl5/2ain5dRhNfr7bJgFDEclnskO1xbblqh2GQ+t
AHQI8fChXzoiJS+/RsHy9JrXPxd4ARl+xqbQbqzwUe0zLLtRWRHFez8JNpveilzu67dtk4DYRrs+
tkzLzFemHMLslAv56s/lEvGvMuoMkJmlWpKSWTMKLeOeqDVospFDCQwWEk1R3trd24ie7lgqcGWh
Jzg3vbHU7njj1smiKPmJs/7cwuQK8YIlrSQdJThzP+Df3H/38mHqdjYU02u9kheGO2pj3zbjX7Ct
BHvuGlaiHvVPI+Mv453M/FJMhkRrPnXgkmj62FrWmhEggU8dRhwOkSPTWvlsUyXxvtiMYruSDAFB
GE/MOtTR7jqIpX33gX4a1CJ0CsdJueDHbGcmtKWaUp5jAjY7iBQNXJPC0iWHxXRTTyL+ombnFGsC
eaYDcUGu3FO2Y/Z+nk23i2Lo6Kpehlm4Lrgz4YGNs/2GV3IeuOSkbRMPBkZQiNd/H7KZvohGjI1D
Bc8z9oNIl2+Ge28Y6TBnhhgKYlJMIXUO1JHvq8Qkjy0WveQiRHEffVlcuhpoMAVzt/vTN7hdX3H5
cNoySdKVD1a9nme8281Ue2pBcTOsZEHJgnQyOWbJreRsb7pYsH2b8YvbdoPI/DwmcMYCF/DVGDEC
dDcOJSOWTxVIPRtbYm14EWVwM+e6bHOktft0OQYvgkY74Bu5ZHLiJC4Phy1sgIuhWT//R/akoYU4
Pd++6xeCjDUkvBvLgufJPkSNjpaxAXaRHQZztGXOTu7nruAB5YzBSSQoJSxoSn0fTiaz+9a02BT4
UPCoJ9fYi4LK+q3fajX4/5ssTfw9REwsuEwPKP5eQLL1M0OAgW0fc+F2u/CYEc4GXXnHCzQ1Hvfz
QCTDSvKauFkSawQKlVMqD0LPfgxZXnu1NyyYfr4uEAYx6mNVHdqi24xC2V9AjExCxOYk50oQHYp6
ZIZZzGUX0f+ZmZReyLymkBIAb9OndF2nFvhjg6KQmznfORSVgTolGB+PQNrXXi11jz4YI0aLWY6L
tzoI8p7tl0/RXNhgo16tjxmNSfBSOAbCBW5Kvg1T2eDyxhdeltGn7jLlVGgNtvZuVUMrtEE/dHf5
dXC4qh5GXDCNO0n+OWcAdyFOqTTenJWY034G8/RV5ul5/v52PoeDqjtnSJkfnD2lCTB73i7GlCOj
wx07B+lDbK4dNJpFjyIeiLL+d2PmO2FqHNMmuXXBjHjnH/PQjKX3zD3GrOjHE9YAobfT4CxI1MYU
hrga5dL8zxpwNLcTtyFGpSJW+OaxVnxIxkB4vKuRdIalOmjSGDpxdX6D3vEFb5KgCNPD/sutGv6r
WDeP3+ysIWTBiB/bxZVrCdewZnSu9adxrw7vzalJWdNDg2UWv3D9gakOhIW2eZHiWnh7ggQBShcz
wWQgRV7WJNnyUibkvJ2emuTOgguZ12jVXLQggZnvnYBI7loZKsb2r0i1BtncV3Ph0SjzSlT6ur2d
M1Gtqr+znnF+3JqUsVvn2KFV1BbIheip8gXia4D/JAX6Ffioi6yF3eDQVfWB9NG2WABXsyx7RRz+
Yvq1EOtDGATFhNkUg4vyon2fmP33Y8L1lwxwLF1yk77b9LZJ3L6LVwDW/fsGPZ28IdhJmlDw4pis
MIYplL+qw9LE/NDynbAS28w0prPg3eNcVnJsGBkM6CLdGCA+1kMrPD3TZku9l/IfSm7vwHDt/L/L
NXlW3vnQvhtnkHBDMAcpHErOEQWnS3wqUKthU+/WysUhcn+YgiPJeF2uCUEyN59MEeAYgpdE3FeL
FlIbaGMiUvuUqrafo4Zf79bqpLqYM8d7JkY24Yyni0Z7NAyuqBzgLSW3ipZ+2wjrK7T7/oRYAPVP
S6dXd5GbdAJw9VKgQpd/PFaqYX9td/Sz9iVkxvkvmdg1RPepmJVWFJ5Vc+cieSxR2gLq7ue56/+4
8eBFqgejGc3BRd0FioOjHIqqKbiCnTqQcs4aWk85hBODz3xC9A3bRw9l6UksZSVnduH/qcFOlWUe
Ecx2KzpGZcxRHGp144Vag61ZZ1WgZnryF1UPS5N77NgHYUmWekL/POHrM4PIH5izxE95arPPLjw2
Bvz87MtTzCHTKB8pOPK30w0gbxP7OyVMJ1y1RJ+eZ4gSJtElL360dD3DhisDFpyEIc8gqABcPJTf
25DGLij3DE6kOvCtcV40MkKKcEmDRvWikd03ctq33N4Re6GC7oU7oSKg5pFr4JjUJ6wvQ38Sv6UN
WuHIpNC3aKdmfr31x09Gs2Sofbkw7KZmU4CY8xUptoWIXI2Q8B03aQ9zRpiXZywb+oC86W6v2P5C
rRenAM7kpLWTshqB25/c9XY5jLZOdsG7zKnW/QjEWHVYYnBZlCXuWiANKr6xygq7ZKEkVBzxkAO6
/sp9TOJF8jQMB2yHAULxinWwjVzEehGz1J1inQHpPEVjS2Tl7hiuIMpyx+koKbJsWahPfRKnUfLn
H4/Dz42H7/9L8MAy7ov5AHCdepGOxBbAi1aV20Z/3uClRTcnzKaUL2nwEGN5p3DMx2Wdrs89ARc4
pSq4yjUgw0+t9frnS31PMyl0En2K/sC6L272S3p42zhtSnoIYp8FMI2oOvuTp2fw8OxSUaYcE7Mj
mVeAzm+nqNuKLAU0Wa4tYAIMwHeFOvX7VgDfJCX4uN/cQPfnsa+OnzgPQ4rbGIhe5sODszye+FyZ
YRxOx0/Mp/tEsp7MA4xRhcJ96lRt2gzfQPX/LZeH+TzgTUxhkCfO583TzbIvj8NMePtun29pIrEO
DRECm97tufIRpH/Q8iRWrJa4Vdsiu/kxWRjQhloYj61JCYfa2HRw26B2o4hSCJoqpsd50/KR8g92
huo/9GwBMuOJ5w48xxH+6Ice3KNKLsbLsmR8NCrnVgGxMQc8yrgIzSeDEmN5IC2pVrGFEmlSeOe/
ndH28mcVDNKbUGS9FR6fjxnCB+ybw+BRy6SvDZw1uFsYZeFWcaq5yZ8xmxq7WEuN9fRxRO+CZBQ8
D0iBpSnKrlozY+xWj+FGywl/ycu8TWwpjltn8CRC/hmxGFLPSD3mf+DLFmmBAIkL7/fY5tJTKNSm
S9Lx2uNCOOKS+Isf3fcLDTJbFIINZE/j0lpgr7JfntgAVsFLeL52B6pYPDS/d0ZMoeYf4+I+NqBG
uEC4ymtnjJ7usIqn9D3LRuQJ1ms6EhzNW32TVxoDkM4qT1W/ET69B3g4GMHTcrKcBMiZw0PewhG+
uyuz+4tPCbCjvgSO1R37s5/A0WdvnHJv2Ev2F4uWojLb95ySsAHcmo/aAh/ZV86swW6KvO8PS5RU
IdJE2Lq/+DVOPWZ9HRGJxL4xpK/IbswesKuiuSIZn9/fsdfz4jEbPTH85E8ytp6V65bbkZJIQyGw
RjDG6I3qhei35fWVyilyEQHlUBsgJrkGlC4DIohOx9mNrEbDQZW9DvEa+2oQKIdAZYEaxIhPcHf4
3g/vLGA26CpuRDxs29qGKJn/jfeH3oBRBdDXwbPUOKzxjTKCvAElpy4AOQmx7ECrE0IMUgjPyOfx
7zzrdt2/muy4Skx6O6pvGwwm67Zd/AgPbEcwp4gCGxjN2ErFNAP8vm48Nn0NE5GViIj8mIe5rzxD
iOrmsovcpCuJnCSUwnHB0PG32SSfA6QUAuDemvgDsp4xRBGlXSIaZO+rZkOMKEgIrFCZodQjoav/
VVXlf05kM8dTCT6VRrlKwBksv4GslUJXecO6zcwpnlbWgwKuicYkRzuzkDrIc7mrz0C2ZsWsGl74
npy7d0VumvFolYV1LqILw1Npoz5zikZCt48qjTBaPvJ2Chu3iRKoymbJy76BUT3ejDivGtLfPQm/
3e5BaVWjWndwFCM3pmlu26STiFmaUq/DHhRqOW2PpOfC7qFVbqr7Idf6yskj1PQCvVNL4LQdImqP
954LB1nzzcQ3aV4nGuTmpKUnB8X86VuKtCWjWyMyj6YOM/EMcwZ8asvLe7MsUBDzwE8Ceo+d+fxJ
DdRgAJ34s5WqZ3/gD9T46XnVfF0bV1bzj4Yy/qe0AJ/0NQdMCVdVLEl5e7OUuZHCuTVdd0RCvn4i
bo9a1IsjnXDlAOd4GN+8WXtRe2M6Nnu1OIVR4/tdwOEnD1YG6sJuNHFboWPmlW/Dv+f0afS64tT0
Xtd/VcfzBUss5ZDEFr713iGne25lvBrP1dX52eZcDYnnNe0j8pHRg9lzPffYn2RdZE4VvIgcoNi9
Ir3GYixRIkUp1UHxL/zy/9Kfn7XO9jW2NZ1S1EJ/E6+8MN0EZ/NHaldtusWCc107FMVtPunPKONp
XrWrS1nxpLWjKQNT3G1KRw7Y2U0AbYWiCoKbi8vWrUyUMgebHDFytFSuuABzyVF5lNWhorQ0x28W
KeQG0s6oXNjB/umEO8MmwPi9QOIek3XnXfx0H0MKj4lffruGVzoMjEV1ZNw7BFgDZkwt9KA8BMqY
6MbPgx2t8cYoz8I29yvI2OgdUnYxDrE9Ia6GGmzyay96CjmxyNRvQGevCjX9CIoDPcaBzsxC6BqU
FVNmhdoFHUNtbHDUgq2Tk5K3a6aXQwxd5zvOfBGpxj4B9uq9r12eHFUN7hnn9OixIH6FOmpTwpp4
e9h6ghs/2icTKVK9a741KFnO+vGTRx6Y+i7ptEi4tSOMnMFZTfCayO3svlMwS22jq1dKp0yWwyMm
WNecAIToAdwbgPPFD1cwCxaONhXCWFvBACPLiBDHMDYYjNSXYum1fN7CCQt2BFqnMC76r5CAF7XC
BshUPt2maz2o/IZWGb7tTNScfxoQukVXqZ8fo41/lFCqSMT9T3lyxmbiWGMGiPxeKO97AR+VzgHd
tYvk9WBUZOdnUaBUOZiLDCMQppxI7NcqSs1uwox0DoxGafylkDWMEHyWBUzcNbBn/JDy8t5HU550
xqAMgqx9P1Un1GImk8aeHLSqPUZyEOWIzPlN75ds0al/G9yd9479WSS6ktO0XKnYXqwL1LNz+KZy
cLR90v5UC0OkCqBWeQIBQYfpGwjXzz6Fooo55X0r8YCSZMfvGWwW9pG9sNY4znGOt6lWxmdvuNzk
C49W0yIFGbBvemud5TrDKwrHarctMR/6jWmSFuZfROEOoysh9JAcmZKGeqxOhgvwJNXZGCfDzWAX
8vrEGA5Qz+WZiZXvIoCnz20gjyWG35cTlcrnJtd8HBkEnVVg1mJatLQPMXtV6eUa5VxwCzWJZX22
gs9aBXiS5gpyktNe16FjEu2yUyCo2gkF2OCIn5HOJUQ8u2fbX0kpfihrtMrwdPtYMsIhtkztEpKW
hdNeLlPqG2ySxJtrw3UDyuEF1vXbc6bW3Gx9XX2szBbeYeWNOlHAVvtlU+RZEgI3nshXjBpHGyb9
8m4DzpIDYSPkbjWrCyin5DAhkBv7gIZmYtPFLQbjx1MYZUQ7bK0JI2mIZCyL8x+XAbXOPr98CnuC
lft3n8JbACTZi+3rdZ14C6XEi1o90L2J5Z7wj5Bm+EnT7rD++3Gxu9Z/paog43uMil7TZpmURCeT
O0vMBi3TqDFQ72ip7Cbe4G0RsYl1SSMliQjBQeX6M1v2G0i5IR/g9gEsn8XadwIyp/COPD9adYUD
aDvbYhOyphklPeSGdoqO0u+pGV27PvFGe4xWkhvzFgY/HEjjr2NfubYjhz/tQKiKgLdsxmhO7dWs
LgFD0khfVOMRHBpbZaBq4vHUiSukEhrOoVl4IpvNrrCmFsjd0Q866qu1PUv2k9w9DfldZfQhxxmg
/BTmGCRjk6dbEtnGhCGDNRa1vv3fLnPeX+jboo21jFRjQ3XTJkVyaDCTAJ8gcUMnHBusmJC+Evp9
BTsN4p1y8FNzIuvsImWLjzECvLNrEYJdi/UOzA/wjk96WE2ZHHrsedaoV6wqivBqZ24qsp3ktEXg
xEBMfUVZKiu4kJ66+Bq2GZZwuZBGy3TlYBbjLVNOXQ0hKs8gX4rlP9bTwN/xE0N1RXdBhp5Vehfr
u0ScHjZ3apcsvfYZt8UniljHPytwACPuoEq9gj5k2Z4hk267OUmXXAHFczXjIhiHUR4W8mxNGtqh
tsIykgYb0VXyGS9aZKnFylwuiI+BZ6n+BP8f8tDwlrpFa3QuSe2uomjm3ixr0aI/D5G/TEFb0uU8
ufgDGrQLSiW8wsWu/ROV/1md94b7ef9BwYVoaFkrA5Fpxph7jWmjAcXDuqslHnjthawQFEUaOLII
eekhxQyRXDCOykxnV0GszUQRQo9O/esi+FvmBDeq7Z5BJdo96K4vO0wztWiwGp4LREYITyub6ZjU
9gMsWOXKFZOOZCXpt8Qltg4mXl2krWzEugDO9gyBNu8mvrE/EWW7C1ImKnrf6fSHP613PouO7Do6
SxP+b0Y7TzboDWyubhwiVLt4dL5AgxGMXjrnaGKskkyHLqazN3y4yQIWmW9OE6F8kfLy1DJSBra4
xMBbKv3rJ0mOUHUyQrsanI22t+Vg5rnwyh8Pm9pDaaEpSCv/9eYDW2y69ywHCMiHdjN6pI+0dhuu
1wEknJCmDshJKAOB6ToRifO8X8GbLgYnOICOzdmsI0sWzCftdCOoSlN3QqVm4QbNv8qABCrWlgC5
bTxgoWhvE3ZG+TNC6KG8RMfy62Gczwnss1pqzAYcf78bwDQFCwHYziDIeDH5ZY0bBYnkqIaC/MZ5
ijSPqlIAl2GGFY6v9Cn7Ei0yArBn86VbZvmrsC8NIqoJlRpTDomLTXoeSgjQ7EpM91VP9finAmgt
e0QtISWCFF06G+5axSWB9Lru5vur/4TI/nL3yOqBp9x98NT83ncDDiV0Nhf4lB9o+P/fRQO/m7/D
iVeGe1+xjPNZGDRAGLMAbcoTFXCqMDFppyYopDQ7wzJyEKpCHf/tdtuTLuJHsRIV8TgMdcHesVM5
+JMnzFqgNbxXNkK9VxU/3c25FATe80QcpJvAqaSawRzljpcEwYIoaoLqFrvhutI56Q3neR+3iKOD
GILHW/8+AU/DpT42YtV3GR3gsqK2XrYb2DVElghT12fn8JcuyeBgDLbGa3wZXPMkWiAl8EkqevoR
VhXbar4KVLFDPTYcvT7/BLxIGAqmDRLoQMJol845zN/BQReD1+sXQvUoU2voDvgPszuAb2A8a5BH
t2XK+W/dSQdGh3MDGy5NpnKNqmyiSXOhVGV4NtQO3APKgjzqgne3KkV8N1oxXicLFsejsUB+iRZb
RKM0jwxFReS47X4t0I8zwrHloVEo0ZPvzc88GwMBI/l2kRUeuovKeGBSkZNPZi5LS/bhZ2QIaqwd
VWi8WRG8XzngUj0jDZyk6mW+yMMJ8h501IYJ14ZYGlKOW62qbSHrVTnE7w5I/B3NnaMilD5FA636
1n1KH+83vQOp08/4veLUH5yxMTQ1CLZFBPCdajANue8VGrI/jzvHvYaPtoFz/y+0RBmyoeDgc4Gh
c4yxrbpj6g0iM0+jjMtInNcmJX/BfHSpAy8lglYwcjprBgi124Hl6ADaWwgDtmkao9u05BccdKtb
Yz3adaTIrGmcoO/4DGTN+aLedR6CmPvlCTNoiyKkVzJLt0bkm/MXA5hFuJmQ6JYF1z+MO+OnMUTR
d2mV3ex6oNCHc2WaKa5xQlZbj7k9Llm9HmdHrRbm9QWcZHm7a7VYJ9ucnCa9nNWvzfyswvOVccXQ
7iuMxyRL9p8NYHtkeijA5W/2DYpVR3xPIW3cZ+uhzixWPqtVUOPyytR27jaJXBFu2ctCZj5/nxj9
UWsM5jS+d4MGvaLgmpx+l/+JbDrewPTv+HllYj1t9s0o/5iDbap1Zoelb5MwMfC42auiUwbuz8WX
qjaijz4PsyxSvrezcxyi92666HcaKSZcnf3SEbGaxcyPdXljkCv8ZV7dUZWYZTe9wGVoWGCsJufp
1JOhb8pshg22/M36ZBB1G7XwdRBBqIQ8Fd589xjeSPF8oMSdk/9NtIr7Rq/N1bftbfFlBMNeqojs
01V/XbgkRk92s/UpNJvinm+5Pm0jOpkOn78Fia9S95boR+r0kYkcRwH6CQLh+9VwWkGh+PZzE13z
TllF4LcJBIU2mTtdO61EqITiARs4dWd8EqJXXEqTUmqlcoz47AuHy0cUuLCqXKHtmnbTV0vjDvzZ
bXG3VoZZOYIBQYQJYWnf+C+UZJHBEErZke7TtxoHlRA/1iI8ArlWqMCldpGLGU4m536Pk2z3st3L
T4cQWROIwo+JyDarLlaVVE1DkMWj5ADjOcnGcFA0LEn6cQW0YoU3gF7V5A4H7+X6dIgH729l+pRN
6hHcbpa5EF5xWX5L1Es+oNXoOxTUiAShhNT3n3FLiQn8GrflgDm9GcxfD2LmmGs8utqEfx3J1PQ0
P8QbzMBxMxVsfMD7FHiFGgsST6NrJNkTLAu8Kc0VS1kEBaYhSwgl1Muk//+iLDDPM9j+GjFScoX4
LBtzytrDK7ANK6Q1APi13roEq3eax3qseFNCe7a8/D1pdYkB9U+k0y14h65/YBkqLIjfVmu8ZWy9
KPWLIBM04s7n/NJv6aBNjJ3es9+CyDKBfU/enZwcvz2yBX3YYcXAjqf6lkSjhkh5kRpi1FntCGnz
Rh0waL+ZjleN4x12MxvJRi/m9057cc8zQXxX7APsTxGYyAGawtPg+duJQmkNthMaAoGLSLqleCR/
eznOwI5+dFAuLVaXm5BCtGikwyCDviBqq0z43SSV29LJ4RmrmnG7nebz7++WjIneffY/sEHPdyjz
NAoosxKxM8+KyIh6p5JQbLl74/sYHPdw2b8qSBLtSqim9N6L841XJBA9iGHLMYs/rcAsF1DBY6eK
avX4sKHcYH06/XzpoK98wlkercRZrYga5Rwi7UQz0mz+/jvv4X59Ua+XfmebxCQr3JVF1QWA/l4e
TosCcGcFRpq5GOlGBvTnwxrvJJIFfJqzchJg+d2MuvakDNzJPrSvVNTD/IEyww1I5ZW3aFa9a+2O
o0uJRWcYRP7zFH9jEXM8jz+tpMsuQZ9cWBf/KjsEKoGzdgNGjjxBv1MWlR3KFjZW7c9PUAqcdKAr
wpL9TTYmK9yRrwY2K8/gcDBBU8q54DMIUqFBy93ML2bvObguV6p1/rUVBF80Hn5IckS4Gv3iu0fA
Kz5LT7QFnk7qQs76TE/EPAASaQiw/J3yU/X7BMBslsYf64guCSIt+AZUwibB9cQlDHcq5xIdyWIp
QPojb2zT7W8LUKpofa64bNyCW8A1mfY02Qoro5bnmXqZNhpWcXkOuTl+xeMdtPKrXqzi/6axQYO1
ugF5FyvkLzgP0bxzYxNv3HbFFjwySxuWcefR5wHP5Ud+B1B9FT/seJVH+jBrQ6n0dy+blkJo4Wan
OcDhiteBedOup1N9QJ6jrz9JPzsmf+dY8SqfyShBJl6ihBGO0CNfjtG1T2xIfaS1YPJKqrB/B/6L
i4IERaGjqqJPl/qS78mg/419KENR4HCf6Z9IUzQWyoH9H3tKERZVzReQ2fsVNHQqpBQSVAwOSfU4
0RRTgMlsFh2IcExUADhXqLVkUDc/AL4E+tzrhdLeDIDgcsIH63/1E57RMWpWHMfjXdv/RLI05RII
DywgHzijvFlYmr6h+XGJMm/QOZ+wNAnMKz9+wNVzPJCK2tfywS8jtZpLKZWx5qSsbRl0iGcbWMwW
aOGHExMarBc5OHhnm6TjgswPHnJR8IGidFYYgG5faOltFoP8t4rgLZ/MuBu6itV2YRjCdoCYy5iK
1TlpLzBO9XR2gC6x5/jYdgQnfo/S6RNbsJQcf+F1+OJ/OaiBrk6ITUnoSar2c0qVKzAKLE2W+iep
eKNNI7JfEMXFnUmz35RYuhfL4mgHv/6I08FWUkMBx6wJCDsosnCkP8m7S4/pnqIUnlOQBDCVM1jO
ueJ5JQ/8EPEWjZ2KQ5eL93x8UWRAUnCMqzblk+NmpsEGBfLAN9sk5OiHdO1ECe148zq+SMCzv+ee
EXIFPQYOy2ziVdYLp9t7QPNp9SZw7BobsveuBQyB0YNIrnJcdX81w2oPOFIB+A7ldVm5eLBcKzra
s1JkdLfd5thGa22ZrzSeuQEuaQdrsj5OijodYggw2qGrwHDypqWrjvvi8IVQcebYm6kft7sv3PZf
QrDN/Lp9eTSYLQlsRfG9YTnajMXluWs+1m+uWOByT8litWUC3rbCEB1W3bea332etS2zuEI/fnfI
e4Fpo1Uw02hrVrlY86QzUymZ4DT2VvOGIQScIe1okZvJ4LEvmtImurZ8BunIGduFdx7Dt91qHWF5
jzxXPIxZ07mu8I8TbQAALcFeCKVAVYbsJ5iXXNqfbMKFAacMQG34aML2iDgmhFxWpwstb0Ima0Oy
bvuUGURkwzSHkIjpCTOEQZMNKKFm0phDcZ6ul6C8mIAi9x2mza0nuzuoF5owo2vnFe8WdRP3jwPY
r+wUEHJmKAYTp4R/TUBpAs8yLhYFsfQBytPl7Ojag8Pwt0Knez7wi3P7Cf/zg25q/GAWPIOUiPjq
xhva15YwR4JdbXp4v4bTnHx0gI4SDdi/kE9Iewxp5iUuTek+Yrc8x/ugU0j7B66flCdPSEN26fNE
LUE1nFKHs0VcXHdm0N0ey+O1qsTPcld2o1GzPgwCo03Du/wJD8JGS6p/1YFQOxv59ve3hppIewr3
RH7zOZioDE8AQdGxPJ/LzxfUwuN+0Vjv7ikHbsXoMlOQWlmVm3FGIHTsH/ZgS57cZjufVK32ea0b
MTVTWL0qHlCMr6TVYh7F1fJ9v5q77QRDDdQRm2Oij50M9XzbNkp82ojFdijKq+AnKnYohDe18i82
TG3ZRdnJ5s1k1Kz1VWSJc1Me47gMIEo7qMgBCwNmbhcJEAIMK8UC/kpz2EMzujigAIv3NZrqPxeW
mW72FjenoS6swlAVxop3CLCDoXxbw0oMkkT0yMwjcaJby1KqKc+mcuy4lHlb6OubL59n/ROurNnt
r9xUP3Ab7cGv0D0hc/UgcJwwsyrQckAVftbQDKOoS81PoVFdMEDfT1/pz67W0ybHHCCf/yjgZ6WW
vD2j5ibQW8NtE+QJsfkd/evkpRfum02t95VRFyj+/yubTTZSbuvCdSjkymvJtLFu3SZ9YE+774/i
jm5KDHB2c2WRYKWxL23OdHmU/csyfXC7ijI4iYvMb8iJ0AxRQKvMLcAlUIzho2Ovu7urIVAmmzL1
4O2n23WhCVTd6KT38W8b2A0K7j4v1phvChQXDqCcFK4gXfI7ztD8PprO3hfYxUGL3ATHMYBijtLY
KspdDwpsw33D5TGNXh8CGVogNrzCe8pRvuGV+lBrr19r3+bvyvwHxHX0OUIqi6Ub1h/4MSSA/3Pd
VRwEmRIwpO9D1wGZQCv/Oa5dDJYKz4z56NaXfneQ5+zvJNCwLs9iFQlD8TCzdBGC/d3dAqfVkngO
2+0fzUEr6KpFGrhKcEUBnYormrDtOLhhoyKvvA5chfkKwjLiKKtn0/SWP41lNE1IxwmNoMVCOkoJ
NOQFpLwa2ypQnFpt17ut+yvczBWgx7eo0ZoVl5BoZsnxAuRiG1YQX7UOQ9nPCKMwq+oWiFg9ndWS
whQV/QXjAEHh88ped/SB3vIFVLEDgwHf3ZdOoSMam2ajMGThw3I3PEJuRe5+E36PZNovu4lVXTTB
/8EdEJAhGCqdrNV+rYGoAV0mc2R5mG7IRoDApMOSD0O2/g2PCtPboKg+bElsYz6Oel+SATS5lS8L
RYsYbwcUOZLvVQV3FlJpjVt2J3TyDjZDk3+sNV8YNWK+iehw/Ljm+8HUTc9+MIWTakXzVkaGboS0
y2e0qfXMK5e029kow67w/TRD7QoL0ADtIm4wXeHXImNjWD1VjFz5/B+gQm3L6B8wDtX4DdFNtP2G
87z0JdC6HNFOlpr19NMv6WDPDmVCi9dZoBILD7FS9pWFv30G+HP3tfjNDoNJdJtE0F/x9nK4P2EA
bUSxQ6s+sOY2GtiyZ2/urDfY/S0OEY4sJGdmFhpfi5vEL76DNIm5Ds83yBtzfojbVHl+b7TTKStE
g9xwaQkgQXDTUoV+Grq4cb108y8UYaDkUTAcIhT5CypW24Meju7qLFqihjcps/pI3nhwG+J90IT0
rXZflNY+2UYAQoAjZPs0Rka/m1o1ll6um9cQvMLl30FhEzJn6Jb46onZ8Fjl9p6bVkEghB2W/5B4
5TEyjtkqysFEtpelYgr11xMMxZLdTquaJkILI8PGMS9hFTxlRklGFGRiKzzVnqczTpoQpfhW+uIP
sIkd+CEHnbQbu0jGtJl5l3KfUFLhXJEWs1zvGZR1pkoPeju49aFDfAKEOrochUhU8m8aWc6vkRSR
OJVqZ1o2DeUIK+MQowyok3pvd4wfJicugvvoBiXYHINxmqWh5V+iAgHO9BAKXjhXT5SmMYhzLurB
VMcqNJN104wd7bq9su3rtqE+3tLbgDX4OKoLrs6YIffM661VllDhccEqtMev1jDa5Fy/dKkqsoXF
Z/xSCvWjllYIJzydPJIP2IkjE62ggl7YpjG4jPXvpceubZ7vvjBqznycpdutYVOb7awcd9OaTdZR
VEcErs59idTNzeOfSyGECfp9ECJFj4cE3CslQk9a85o8pwPjSigju/O1vZPRetHwy5snPywr9lTv
IMG+poJlBSNNd7wZOwhKPsLcxFwEOCUYSYcAw1m/mp3dLd3U81/UzTRo1Z/hKumF69jxhn7aQa3m
h5/0sHLSTVWxv64I/vSqN/joMPcHSrXGZch0K2utdYl3E5Dd/f1f+K9KiViFVUZ3g2O1PJGeX+Vb
Aetuo6Mpo5yJPCcJD/ezTle88xM5auKWpUAoUIUmmFuXVAq1eEYyG2uuFxG8mcm/P2++Q3BfyPkC
vHo37+7gXdaLxXvTP30ovDqB/XLHd+4mIbPDGNQG9TWrctPGlYQ+iz7DLU6pFXyLjHWzDdzDQmiP
JxCxV/rmDsXMicsstaZWAUuXzeT6nNyXypjhNhIHNLNAExVXHlTDHZmLXORtvqS7bLZ3mQtQNoNZ
H/M2eGDsdduoxr1GQ2MXI6j0ixSQnc6OGKJ+Ct7Qy8PCt0LuWVIB30+ul5OA+r66GijebjWjbLBX
1G+yihgrOQEAAn1JawOIFEEyWqRUhKQpqqc4HCT3wpzFQVBDyXVKg6rJRpDHLBxUOZLaDK5cgdWS
HHDTXCHH4xaTzDsfifK8E6OE0AWJQ4iyjzOOQmDGxDdO+iKt1w7Iao5uHEnTSFu/rqaB3/mw7kw5
QoQrX8vgYhSgkFlU9sNxelcyAeFXeA84wr77kPgSnKBkflTNivBAl8lVVSDppNPe4TShgcjAv4sr
9kCwCs2/A5sExHWFUE9OR0J0wo0xodXtEoHFPT9GkY2ayroNqYpsJX2yxp6DCTK0TUVj+a3HKFWm
9OVlJ8+iivIrFeWDf7VZkNV/utj2kiREvPuzKjqsOx5nK1L/RrZQs6aXT6CxkwktGfWvFvs6+whI
FckCIYNwwhZ3ezwGHHt5g2Z1abjaxL2nshH+oovS3ubbFT4/NZ2H3/9qr2V9qLFisRhlS/YpcUNJ
FKigMyb3+ui0R9vnWlmCO6at4TLsxCdHfC/br8qijEs3s636/fEtMlfx0J7AHwt8XRoTxYdOXVws
25qJgKIIQjwmIYUb1IRBdYs/9CequXCBYSWaYC1WDcoNgbW0cRK2WrzBPdlXFAXyh6Tnzo+AxBy3
bVS1qJ+aWY45soDatYGydbBxWs25vpTfAV6BXWz/dDm2BqfxnLRS2c/QxwXJjEqdaTD8exdetB+O
g5oUDU7yzZyUEoGfnlsG4vqcSb5rZWbm5TRQ/iGwIYBgkMe+gu03Fp5jIK/fSEQ6WdFjQLC06o47
H0iUy7++A9SYE8xWHHKHJwbSXgQchkxPoz/SKNy1LTtGqFBq+enxzpEU5aL3QQmIQMFOqhWAfOgI
rGf5yMj0RokayryvLZTWrtS/V1McTmGk3QCUrIUHDjDeCD7ItD9Kv8fLGPYrvYH4w7mXph3Kh22r
+WFlAaW3qRgWGYUNpz2HD9ac8JthBtEtrv6M/BjOQE0WWkxfwlxKzClcdW9ykEQYJrj2PEB6sE+P
dMMbOcyctlX9mZXxLu5bzuRnlPp2mFnNw/bJa40X/7+HDTJqIH5JP6cPVx1PU6JmDPl9vdcQnHrF
uXEb8QSR7pp3sbN9B/c2VwEpPs96v2gnJFsucw88QIWahpckxR31wdwAQ1/RBxrhfzs+grTQn5Wy
uFMLHqVSkgQAz1oVIZocZ2IbjP89o43k6iOpkfh2QbecC2fD7+ieDzeFbe0jYP4gUoT+EPq40Zv4
4MZ4QlzkTpZWpXS/T9lexCR6g45b/BRfCDhea2Y1h5K4Tl/KJuMuuRX280yKhMlvWRgJdd/lDzIp
KaeoHfTE70LCVnU8QniDA5WcnfSs7WajlhddV3fgTogOcIMKw5+3M3lQeOaZaRmNZHpt675oyWWa
uT+ZPT8dtCpcTuHlsag/chLB4ORz9d3IQPVXXizVcovW84Gu0kUx6r8/6rH9vReSn8ExgTTb8Uzn
tclh9DWq8BGrD7DPwYwTYCr9kF2S9CST9+/N/coyVX2HVOCZwxcEHLThyiGnGFkmgS1dBbikevWS
prXoUNd9iGiu2aqqZlKvEZueQ2FqTNoAfgd3whD/FAzRE4n/nxfiWtjD7xMQVGGPTpu2ja95BB0r
C4b5TlIFaQQ5MyEAQdx+M9xMH1FZSOi0WakfgLqpS+JKz5Y7yR4grsoJQLDPZd/p6FzY0XK0fq3+
uwOe41q3GTktgI7hUV+9ykBGeqza1U75/Lsi9DnaPoTSVI9pE0JsAxIBqtPK35yVT7Wqril/wTMu
3+IAxb1MacdS6AHuzQVt5PeXjpGwU8i2iYrXerxsS6kae6DKHAjxzw8ZpOJ1yMEdgNUo3Ccea0aV
KxQJElIhxSOH1qrgWiOe+uQFJZfUBiSDnPwZ1k0Kg7UsUhB/Zf1VjJr+KCBSPetvwNZ2sMoeBMIC
nWv0CNfsLgjnPktVMyp6urorY8W6Ip4wiGMzBv43k7XWp8ESjEDdpJv7L/BRm2DcBrSE3vFpGISc
kN/EsY/oMY1Gd6ZPemaCaQXBzY+svm/fQQVe0C9nz45uR/wVdCNtSXEleDwNHVLdQi+ax7LcVpRB
FJKnrmIRU3oavDFA6zRSGN/lAUM+3AKmP6klZQ900heAMBuWdBBGa5ctUr8u3tjBvomtWzQFWWK6
s3cgBqOYAbCDHqruydIEYXgytPRH9Jy8CiSzrzpAhy9oDFC35OF/THE2MpaFG5ONnjJv3oawlzDv
Go4m2c/bwubf32ptwoJH3trLTS88eV6u9NNts+3DrrlC3E0pklhZtb1RysZ8OjSXvgcT9Fe7LX+T
VErPceQQk5aHG09fPf935RqrXnJUWAvOUc5PAccUmtizHmFBy/P/z3vRRxIaZMopDLgOtS7pdiC5
8T0CBHJAkI524d+vqPkqJofVZNtMBlRVCNc9f1cQaAvxWNvu+QQo3xpnKITf6hiE871bljXNqjNH
T33/3xR23CLu+9O3L5R3BU7xnWbuB9VLufdFFW6M5OIy+w2N0HRBbcnJ6eZ/cL9YMKeypXOZA2vt
iaig6grAp8oHazZPbdUfg3eBabn27zC3xjxFpcgS4HQy/tWyRvamZ3hPlKWHLmZYHISxk8oqghSX
SbUFXlQdf4AdnYIUbChRFEyYsX8WySvih7sj4MGiYVJzOW0hvenA4WoIgoNTOMm2u+EudKrxsnw5
KAtkVgNdngooqWJ8C7RQt96tlAe8/if0sXNc6jrG9M9m1VTn/37vUEOaISZfOKldhx0XI/AeDa62
3Zl6z4zua49nJfWjrvu0l+2Y/KJGNDB0KT0KdKnt6jRISW5lQ5h6jKM1DTW62I83cCqeSNQlZWDN
DAjSX6Y6089KfwNOy2bKGXU4Qnrdu1h96G83ToYfNp17aVM1mMZxdhmDYVnVWOgHgZgiIPKEhycs
1g6qpZHXy1CBmgn16w+/EP24uZFS4dNnxN0qUXEx9Dw8bf8iuQe6roSWqsRolf6Jf79NvJr1lotr
SLOCg0QgyNGeeDt46/9/iQVFuOWCLXQg3xyYBZzx0DMZnGQTuOuGGoejGfK2FYI1mSmBIi3HPKXh
Joif5UQauGO/EtDDRY7Kdnk4nCeZ54EEnj2IiNn+xdyBgxrWjv3/RY4D43aW0Q5VMV8FziYvnxU/
EkBWXkOxBS1zufh78BHFIjUhuT6MwF/EoGCjA99NZxt+vEPxHyJitWOMdZyO44I0HTi4g6q+Y8CV
MWo1JfqtKvBgH7EHO0PSrZZ7Of5erT9vkt2U+2t77zinxM5ONM5sGO+uBcBZnR5wVbn94qGjM7uP
0HLT43fiz8ouMlqHC7DZvtu5w05t1XUO/nZCMFii5/f1rzhnIf/r8cP8mHPVzwSFRoxLxxu5CSHh
v6C7/Qa+faWQtTeB7nbJHntjiW22SfJg3GjNgj6bhCuKzsr/fcazbop8UFRexqNSBkZIWMZumCyn
lQUpL76Yb53Wo93z94JAxdxEVHyZcXvKW9XNW1biDPTQ9Kxnql4p2yvxJlX6msE2FGsWwzgeM8XQ
LuMVnkIY9scLwtYfcJmeqTp8ditfbJu8rbyi/QHibf8IaodvbF2/RiPtzTBYOUdtEecUyeW/Y0ac
7DpG/HGmRtnwzGAqaK9EF1Pcyk/WATAheYs/2c2ZlvCV7QvoLsRrQ7VdGMdxh0tkPU5rVMtK2cm1
/4WuQYJMLpVgoyOQoorhT9qX0FkmgUgZNwqp38f1IHedatYN7nF0cwdblGRGlCJo1l17bqvb9aid
BBluO2H6cS/Q82H4H6K2lhSOAEwlaI5QUX7U/j3sXCIAiR9DavRPTOT9lOzJREJi8OsAGJltZ8YY
ohXkEgcV2kfry17eb/Rfq6vGbteM4pdVE7Zseyr7qztwoCoCRLbBz4SlUXygVWwqP3S6hZbV5/HH
W9oXl16s2UCkmvDIU4Kqeoruj41jdTuJgTkICMkrF1D7hPJeNHmlH29kQmV67l4rzMqE/zkWm5Qy
mG4DwWFN4OCeXG3aHMU73SZhZI0KN8PWu+vWy2pETuY1GLzX8d9rqcajI900ELloPm5IBghDXxH8
LFCvYCSmmz9WyAo6T+dluUs23jUeKvgl2+UkVIFW8z2l1THFVJOFrScajyxzJdiRjQnA49/WWxj8
LlpZifPVsIsbgeT/R3kGrPQoXFYoFPr6GVSiU0BncIobyQbjVVBYY1HDaewH+47nbOP0baoKaqV1
WNgOjcaTmssKNfc0tO+wXSwBYoM1zLvbfwsXUuavXXgcMhJDPKHV+qUNhulEmvzxQMXaGTKYn75U
JfO3BxRrToWtX8icbHwklmzEo/jTvVczfcvZGDTlyNRiP7LH0PPskHcPNWMjdaTZqLGYTlUitjqo
M1KpDlFWLsy4NRw/Y7TWyr9/y2m0ByzKF5eveHYACxj9+amQ+G+4U09BP2jHHRvrAyQ/vtZrTMUy
AJkdKNKMurMeRvXZNMJM/Yf3MksoRr4wN79WDILQpsfVme1IG3i1wRcKWeBxRNb4/RRyZjQsPBC0
dJI9KPIbxW+UJFE9kBH3mrdWjOyX4FgGsxkTqpTeld5toKL1Tk0xJJEjTqBX01Drsgb8IA6EKMW4
3YpppP3SMlytYewjfXtpXx/OB9UuG8OhO7mXmrBzDzqn4c3/EYe6XYoZNY2aRlSn56K0zlRh1T6G
eYfnTHAtuCcIm2j6UR2LLGh6JDTa4JNaU3oEhjMqGwxDUO8zN9cRbvKDXmJCQf3FbkvvPubXNaob
i+KSJUSIGGf/+DYSHS43ldJW0YDwITV7IZMrXSrXS5OOoGvynwUOru/MIq2jGbXugpToZhd9lKT6
535hTKd9qPcmZkcESkvFgRaFoH7sCWS0aL1826UjNCk5tMFTJB00JPvhOUvDziCssGsbEoaR5ZlV
TAYvwUF+1jbargS2nJSK0UPiKDoeJ5th3odS1oMtVp5BCmGdHoAdsqPKpV0N7b8QgTH60J6NJ91d
IUTwDBeLPkFq1ROK1UxMWK9Wq3nYkoa5fHaPxFzexwKAGXo4UKQWFM/t99kVTVdo9ZkTrd4DTcqp
W7yWcSJM/27WZ4q5ZGdgh3dFyrFqYvGxPj7S7i/jr6Bk99zC92eaPOeXKKeKAJSOS5eDwtI3aLa7
LmVcOyMqkgkN7Y+/cOXuz7GIca2wXJ1cDwycT38GxcwYjf/kohzgWc8CbdMDR1/idZAwpTnSdPb9
/3cOg2IC+6uZmIvgO2CgmA8ks1nozB/HBk5fjpgEKAEkGqNcl7JezSHUirZJDGaGNROPZpQXHrFu
4yL+35LFhS6uQXdWmGxVf866nOgwJXEJOOW+FLZXa3zxeWZWD62/7YzME8fQJfSSk3faNBp4r838
nzOvc4yFEzrK1JFv4bhLbG9EDLa1BsAmgNOKmPVUjmBJFtDtB60k5SZTRRwIXObWLOwPrLEyoqKD
ARiKSP4kILKSaeNsJCNR330BJZrT2QBVe6oRkbm+930YXWNVCKzldK33ei4hUKlC6WbvXR0YJ5Tj
VI77Gr+5Aln8UdId0Nh6ZikG9AdcKrq21f2qtj9cylMte6eQFgQBd6kY6UbiPY3wovrnTuqvwPFh
HV87LWp2eyql3z94Ek50PHMwkA1rGvoMs9rTB9oioq5AO2FAg7zgQPR5DoTClBz7jsgovnzw58Rl
goqwJLHp6v2xQD9w+GXomlrvMFrUS8r7ZXT+0Z9WJ1d0CKzTceUa4EVGsLobo6qnPt3kr7AoZGh3
NWVoqYQPP1/1h1L4tQJEFTfWKIOdMcz9mxg+heK+/YhYd1G3OIWypH2rVJx2n+BYMEVZDHgkD1yr
bALEQiTATdGfiJAopI+mj/UlwQkiA+OElJhAzj4G+/Pk+I+xDlBQ7N3X43qQ0GeSOJJ3gwFko+lB
Vuin+yUVoKbLOBm4h1P1cBhAnKOUXuRieyV1Yu6P/0mhAm1mE0ISt4Kc5beyVe/kEr/AggiJrK9C
j+ktLxvaCZ9IvZh4QHJ0lWhkF2PeE1flkFJkVRnlfTYIAuKxW0gXOOaYl7+OcwzZJBp7ED6CVxsp
awSMN15yOh5iilNCN37ojyutkraIPF4q2SlIUyVctyULfDIwFP5pU7yssbuJZFf6JT0bRfC9IVkx
29rmzxuLcN3BmjXNE/HVO+V6JOgPbg3Db2izZUTacBe0So+0zqLcFUkD5eK0TAYRh/jwUhoWgeFj
7gKo/bygqS+nEo8ntBS2COcBUp+wyRd4YvW0oVgcMxVL0Y8GRpbDRJtBSWNqNK5qjaZ8rStvNzgA
to3WG/glBtwKVQrFvCshohPoapHw66vBh8yOJqavvGVyqmVLwT+TDVMp9lMrm2AcFAFucA+MaXe9
4VJhVXDqRGlDAFle7s/5jabCtPUPhrCDEZ6zhwTZBOvei8Hr3QTNfgkpXyyCxmEJCcz4NQmOlhtx
3PHlyQ3NkxL3dzQ90n9TN84sjXxG9nuJkUelsxJTraK4etH0UCrsipmLajc30i4Q4OVzGkBlSQX0
atdWI+0ZmQRuESXrZqxQ1wsSpNOoPvIFQ30xJJPlPJwkHLYmopF2MQQL2kN6iD8yCuyUzJ0KAAqz
odNNFsxJk1bN2IuAswI7TCmsiYfWTKYSmseF6GW3s6gfgn6zDsMRDyuI08CQBiso+c22ExvaKDDV
RaewheVpyhRw8N//JAssk6ok0WWffgN0YQ2SmQ0pYec0tesq7c7G6WIJxVxiDqLF0qFDHh82DWXe
Tv5hIwtHNrDR6AYE/R1ubmAz60Bv1U8F9aX5WhqbwnhhesnTV8nOtakkJ9rgtqmrVBir06jUhCkX
YDZLyIYEX8rQzXhG51J1ho8XfyWlg29e2AMcXFMgoWXe+ag0kWKjUe4FssHqBssZhVxPeQ7Fqzxn
ki23WPA8HXmVdfb4hryvO/Jp6kmbdCuA4uI7mN6QqaPwDSQnGFg+UpbTnSH8Ly3yJrrX5EXHOnPC
KoUSlpQRHXp40DgZEcZa7wFfanAttS0AqE/9qkagJ93uFfBNh2O0hlrg8IVO1TasYomIzRUf0J0f
1biafmcBsHDxoyEznQ7P9PyGABgcIrOSTl2mVHaNrTNMKGUsvTZ44w/50wr/XMqItYRxjjdi7om2
iQ74U6acwMytEhsM32kX/Vi+qMA19h0v8pE8KMzmwdTCuSTr5Tb2QBzTJr/Vvz/MzqjLX38rTcAF
TzudHXvjx6Czso9PdWYdmW1/QbJJDf8SqeCiXQdJJI0K41sX3rnHmPv+kDT2XYD3aT8cdnmBin1P
40W7SKARozwhUZBeWHDgj9811cj7FHODN/6jlHslqG0ryh8xi9tOHNh99d5aEZkVzk1AJwXUNn+e
A/8DFF68tz1Ef4VGza4Q/BA+Wi985HaVHHglPcEI9VI19QNRc3pwL8oEcmYbQ16TzRXIK5gE5NR4
h40ozKIQ/+Vi3lpaixDZvHJT5tRm5cmt0b8tYboCDxv/3NoiZC0Obp7NOsa4N4lhTW6B5YXCKA7d
MqXJSsBXhDY8wxlEofBpv3oqkgs3G3+CSKSQiewm8yVeV12eaQPWGyTo+s/hJX9Z8uyiP9TwDPM3
OEH5NBLCsEElVxrUEDFp8yIqwrddDlf8eyQs4lklcbEwDf92sFbb7Cpuh2vSLA5OhBJiFYEPQ3fg
jc5XeAiIeA+KXuYjY38+7xyTi0b7SU850JJTMDXz7wxZCKL7I2z5ZnfmJTzpElGgWRjKzLBw6G6e
VPxHG0b54tHOxz6agBc/bh8KA+lbDC5ox+HPB0lAO5RdpeOICefCgo2WWrL0go8WDwKXpH+v4s9J
XUCgQdiRZVNSFIeuyIiVxOkqdbe0HEfLhJleG2Q0w8ELFHTNljhtd61YLTdtH8eEGEgiD8YRBBV7
w97zu6xF5aC3aDNFqn81AUV4bmcHOVgIIqjFlRBiwKYL71F76iQ6H+3kFrKpmMFcY63vthEVxuVI
8xRbpOYq0Vb1uI76WSbzce1y40pE10/cUmaZ9KuKo+hjMbRCdljWD5PopY8ibdMxH2YuZAh/2bWL
w7VZkTBoXP26jQzXdQqZC0z4iJl+NUI9qkueiLHC30t82OFBrn0SNFVkdyLcdDzjsn/hTWexEUj7
0ixvKR5U1BLWi7Ygg7dc4l6o62WKBz7gpjYij97PytRuWOl42N1y5okOsEZWhGBqwZpxPEtnm+3L
FSA0GmeWl8jgOejyx5NiungWIjqW8CZiYexOGnlhOULO+fV2Mjx4qxC4DAaNehFn0mARyCX/MyLG
oT0A0mFEENdGeiC240aZGkfDPzH5iUNo9nHvMYffyuPCiht423Jzppi/sDYmfqswrknPkaHATa5I
TeXO7IAkkcKRHDijSHXr0H1sulnSxM6shuLjx0IfxAe2PT0P+WkBan1kZe+bb0THnBT4Thqi4Zs7
ye88O+CkPwdsoAz6WnzDXEPHzKk35C04rNMiOcQaDy61WsJ6GGVHcBqGPSrZyIe9oq4d6tqwiFz0
zOOIRyjZTgUkArp8jlKnsqrTL3uZScco34W/HYdUHwC7x6pz+/NajI8CV9+HOW7BLBLsR3Pwvn9b
KvH93ljhB9LxgGe7zaPbn7RolwRb1kuiCA5PFXc/phzgxR7J0/I6b1Zsd9QrgWM2to30TGNMb6bW
/XV+dFQ3aWOHTeE8j0SFwR5NYN0qqsMIwd+5MPYpQqNhttqTewQHCWvaJh65yOMLTZsMcgSNdl9s
pU0QfHdNvYzeCSfCOJmF29fzpMDYCLwfiXbSjM4PFkxuspDl5uxcUyQiKeIN5yDZHrXtxPTTDixh
z6Vygs0s0nURM1jtlPqQMTxYVWjUjGq0pVyOrKrZB01GYs2sFubBxD+a5H4HCKyDS7nGQgLw1ew0
Gq8sOGtmp+RqBBlFB6K8i2XNq1jKxsW2jxOQb3We1ETNzLTqaeUJ7pL/jg9RpWzxypzz5bWZwYAg
NDOlFRx585kvhQbrDHANyMCVl1BkUFzr1mcOzzd8yGC7TjwFBQpahp67P8drsAJDG/tdVoiIsqbM
KzFsxcmJeybjvQmwarJdLU6NSqSLnWkgKXpc9t6h3WAB4WGU8GANAhOqmzu7Dfm2K/tT3G+L5H8d
7q5TvT5LYNUMN/Zi6lCgz49qW6jjVVLzQ29L+WTt4ycZ5n4IksekMMc07l5YM/naR8Xz2Gauq4q1
YO5mzROS34uLuyD83C9flcHYF8cKbmKZ97BQ7DoiTbwOpk2uD+20NGD4hgq1Cs4g1FLCNAXCQDN1
K4Fq201Uh1IaltEiZT0zRjP+Dl3SRrxOzN+qq9OhJ4ysgIZdgrGV56p343bSzC8O3sjsaz5UTZX3
+IBR9NUSlzTknb9+YjQi0PJ7Cc+lA/1428aaE5w9YnyY2kOP7Pa5iz29j1axUIyLcNt0Eu9ewE/D
Kta79aNyRVOFPxJMMILpweIHXQ+YKFzhjstXwIO6AsjvIuNUvGw50Ju/FLGDnaffN7NFo0MzIu+G
bjC7y3dMzy0P9XHHYOLPwIj/EjAA+soKcmasmVGB31OeJWlR+FVfHBMkp2aVCbCNxc9jSJkrGFxf
NvQwuRnB0NG9HaxphO7UpFXBLSkNOf9nY/jmcLEHrxnrVvGNNHC0dhMJ2eyCfoDgOKl2TZtAuHGP
/ljRNl0xiHmcCN/NdaIAJ1XOodcSeE5554HQpF4pcrN5KbULb2YAxPZTkJaSRggzWWjfrwYl8ZAN
mD1FbjGj5AHRA0FscNRNHn8uJNfPDRqQuJ6hEgYgm1Y7j1rRiPkibU6VIeC+KX8usPbLajeJTLo1
f+FVzDlHrCNFr/Ie6qOuvoyOrgZroCLVKPRFRDQr+L7hzgoBMWOVACjyRA4FWyg42iCejG83QfTA
V2jovjQq7jhNV1J9gv4/zu8SQ8Q+CA9e7AJkFjNCtJSjn05yJJYx0PuOO+q2Z5wU80t+cuwZJuDh
J+2U4Wl/+fe+QVoLwZ6ZIzNz8WQKJkNSM2DdXEzLhKK7h9r9oUIn6uy13pr9xSIklwHpMK8oMEsS
eAIFRtKqMZTlL/VAhvgMe1eJ9n6rYUiNHn6+QmEsXBUuyOVwIsjBRRR2NRIMdkHVIO6eyTQ0Cpju
rFk3wyAoweNSRGnvmlUgL5M3Cm6AVhwB5t6DYmGfIF+iCN3ndJ6YjnMr5i9DYbuHQNHdv30iFIgD
hgCKO0i22r/eJQLDMAi04SASrovqUt7w2/iR/1prInj8r/8ygZCjU49Q/4d7kDa+VOHA9RfD7wpk
HIGn7DOqto96Yqtn/HEMKDnQw+e14t8PLmtD0puygBCf6qxFylbpZ6Lb6XvTKHSUItnfGKGeuSHH
5h6Z2uZGjE/PFSPjRhgT38zA0SsjHz1kpgj/qzaIDzGm1/8Vd7TZBWsoRAkbP6tthNKhcn4+k/zc
0OxU9islCoMqLzExGBXpoyXbaZ2mPrfObWbNTaKbswF9mmqifDfykZ4+TL4+AwQE6v0pAmElyPWU
u9XJyLNZWMjD2PkOW/GeEecr8975+ilFOHBDzMhApnFvYyPQLDdSbKR1Jhte/36CP0pdpm0lisPT
I7B0+dT/8GW5BQM3aZIlNZA/mL60U+2JkNDd2nf+QEDeVczcWtxzrwL0YjOokAePti9yo7vwJ4GB
PCnXfsgVfWhxZB8MMU0XhHs9FnqGyZNPuppSGRi1mKAsT/mhY1Qc7Ys8AEnmUwr8znYMZ1lL0Ltp
7EP0lxkdqzuagQtdnORGFQp/sqjUaP8TSMwDdEiEIp9ANrB86bg5L5gN0vFjpWaMOvwvTBh1NdWl
QWboz+P9W1gtpGJvUJ+Nj7iHIpC4ieaGxokKaxcdo0aMVhn2gDvIY1rUyQrjaiOPJfk7RkAaCrV8
1pXHXuwX/7gpVduFd7liIjBKFvW89TUbzZ7JbVLAd2+1LaJG+3eHzpo6xJ5I4Zx7lAk5ks4s+hhO
XU3GCnbksHV/L2FeNWUvpdlN3m+s/Y5/4bzbLb161kGH0UkZuNrTL5ZE4v6HzFJLC5cMC68igNSv
JXtgBPa3lidFMPVrG46+UxcP/TCQryxJaApY3yf5/tKczXMj/lk1genAjr/6voFyKVvWGhpv+alc
Iwq7lhdIbLr5RpN6UnCqxASgub/fTMLXkB8Dfby0DKcTJoloDUfhPialq+4EqyAE+mKOimOWdxja
+b5SYxm6z94iM4Zz78sPrCZAosA99Uv6lSzxpg2DVnZ7scYtO+qwn7qKjy1uSXB4YORl3jPIJLC5
fa5jx6WSbtoixqn3irZ7T0s+G84UXZw2OufZwdAPA+KSslkt8uUNIGVguOzuMYkZuTYr+Sno/LlR
pEg265RUMnLuEbzbw7OpcqlDZ85922ufzpWHbCzBqDOBdnPAvLD1ua5fnaWy0qdqR/C5FxqroEgC
YcL+/F5vRAcBtrvkhJWgTDFDykErKrWg1hHZ5bRtFzu4ITyqA1TRJcDG10IVGES9hyDae28fojCS
z5nIPih8uK4dtv2YfMzypGNgbL31sU8H/8sFXIM/YjlGlApgZgOlSHH0B4eqYHhBN+ZfGcbIMaQU
Y6j1+TJFqdKe23nIabl3tfTgv+4VmYi6OfOZvjskOKnJSyUdg4Yga5ko/V/dEnBSzSiimb9SBMRR
yQiJO8Q5hfSGflCuM3iOKXjczvpIXHgfkrIN5dhwW4HYEwqWVTa91de9pdNcQ+bZ5DNqaCvP947B
jUrILvd4TSA6uMIHVcZWMrM8DKbMcUeHMoecPZyVh41e1245JPpDeYhisOGVUAFicU/rotEefOV+
S65OnIP2hTBRykouMjiIYdytA+XEDA7iDCuefOrq80E++uUA1NrAv7MweoPFDGMyy6tQm8acki/0
yFPhhTNeuvMOtIDc0fftx0GaUvdPABBpz5R1fwTI62koMI/azd2PUy4OVfEd8Q+gVMc4CtNdoJUJ
m76T880dr+Gi2W+9TWxGRS10D4Wh62rcGVoqq9L5r3MbGVgYTQ6YdO0u6R9bRb15OM1Ucn53w3S4
V9v5Fq6lypYHt7mlqNPv1TFRkJ/mzx4i9fB3Np8nZEpRyH0WZAuh/VipBOs50SMZeD/8dpyFBhjp
rDgRlV5/g6l/f8/HOBlEw2agaw1mXsMSxiOYGcBp3ry6Z+7CE5mOs72joYxLbNaA+lh5p4mCNkdw
1toGSTpJZHkZZAxxG9BBmABLYyIl5kYBZku5yBdDStQRdJ+Ty6wFsNi+xqC8vSIkYMdPICBvxsqK
SE7ycGpYQWrBFeh+Il187BZv9Z5ZV4Qu1RPoeb9FKa3aHPZFJZLAmSk35MOdQuV10IeTCq+dfAOp
hloUVDlq73yweRm6qSH1ozxNqKK3HD3a0jSdwmcIQnJtjRUTOeEADLHXnF+0ZjT529rO5zBM4Qdq
UHO7dAUQU9eb0geuVyLP0+FqUopQ/pnVOEPnF99ap4OsqL2DM/K6RlpBwt7/FGEzl09YdeG9oTRf
jKdWzombTCYcGmvoMkq+JIit7PDQjKsU4xGbCMPXyYejuHtgF1PbdeCIqBvPsbxAu2J+iDm16k/O
pLZUEUxOBrLWRaVtV6wgaxveGJNhV+7VQR4Q1tpVnmflrq4orGKogQtI05wROxCW1992bPo+mz9d
rjAnbarXGkT30Orxe5+hMO3dukqvvOrfgXlSd+3l73czU1TXHz11Rcl+l69+9221nk6hGPe4qJGX
UCzjZZu51XqEUeWOgmYvlnEwArZMSw6cOOYGvPCg2WVIKs45Ib7cusxSzY7apxbT9YfsFcOveWVz
RaOzR+MoD2e/m2TMER5rVLhsQuhjrAfrlDInAubX++ndpe/U1tcKgyk=
`pragma protect end_protected
