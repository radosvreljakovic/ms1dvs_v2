// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
KCaSb52IN42NTD9rWNLc0MA3VM6aR4E4IjcsjhnFulyi0OcKdvtSsUdH1Wdva90yKLGEPx+aNZ/y
zTmZfWmcRwXml1eez/9uGz6g2eDjPOZnN8611MkoFl1h4BtDy1HLwmKLLtUo+siPv1qwMYh6U47e
kJcyFJteFnOftkx01b4vnpZkNMDtmC8O7E4G1hAVWBcFeIE5m4B9RW8NI7rBre9bY+tvTGu23ion
YmNGCLNod+2lquEH8pvOuhqxfrHneu+JBrdPz98CkF3i5MNNFXap4oA9lfnmQdhJ5yz29rTCyzk4
ekGGD5Pz7YVZdurihmMSUqCHcYKmZ0Cuer1IMA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8dCTnLvkiNVgChptjz5mQ0eZP3mi4RWpIf7fgO+Qp5DAa/WfZjF95Axq6v6KQI0KCk2zVkuZGfP5
wtxiwfNbk4tiwl77Zhe18GBJCZJFY66dJiKHLxPJCQF4SUdMtgcK8kMo0hZY9WhLQF6v8gzqpcVF
3p861uzxdkcBy0q0tGX4pw7KI1t7A6bTogq1qPQ+CTPXwtlLON32pQerxNM9d7VpMpnoHmb5cZPM
100TmAgc4WT9fA/R9lAvrOZRrFR0TOAl4O9VxMJ8/M9qwZgg0FFuRWqVcHEDR7+5i8cDWtvwcnAI
t+9UWHYu5H79CsdThTtPZOe1rHbk+/+aJUcUFSO7ll02GhWvR0EuNcs4Wr6bB6iAxkPglhCVOs6A
5caTw8hjdbQPmtCc3nDjJL8Obmp0fSgIi0l0UCBIeuO0porAEcUUU5LPwZrGlCN23U+xgDEsbpB+
fiqUWYcUXZA7G71IGgNvfhzOcsMzenVB1vAsVdZ7msZi3zuAv0tKczHdxznPY/HYqgxrybM3uJFS
HDcW0m/H9yHbJIqtQ6HykS2sMPup6bx5KixcPa/RccpZogaYAwnf5wKhnCtuxYy23S6rsbdUzEOn
KdQB5KSY3KeL2MgBcc0qaYFGAQFkgkXJwu9/yioaUvqW2F1E1h4jZixlWllUjf+kMMALfb6ck1S0
K65tYstAion+H1sLwzuMNzv055l5W66B9jSvAY/byeS6I/uWzzi/ejWR4nWy5eKQru6OlOgVr/8N
cbfKl7y+PCbHehyS9i43cIS+NaTqR+0LQGNTxdCprgrIspPqoEHRoQt9JmMCaCz5vaRb73oTaMkB
xep35V/KrCO0gTtGgXcmAnbyGI3KzateP9MEULhva7drJY7aLwtjcXBbqMsTdTqsRhO2WkvgRLss
1sqZgwitPKUU1T838Fj1kexAbUKWXBW6//a8InUDafJJw2NOXoN1IZdmPcrbE2tP10gc7xJE8dX6
mIcJ2vUg0eOOLF8z9VmLpWQ70D8RaLmYAHAr6hJ6H0+P6J9EiRh9iO9Gxysb4D8skckvt6KEO4oU
ZVfkGCAMZlivXiu09l6Ifi73yeA9xARnyjXiyIb23Did6HMcduEsGXNvXe8jgtN3iAQDcxjMgujs
M4zXwRlqNP47JzODek7Dpnm0S1wK48MevBbkYafwuLvWnAqNxx+cCX66KEv9iWGTIUS+pNPC0Don
Mmo2BtLXFus0F8p0ZNLO+Ulxs1v1FAH8Gw90LmjvWyHJAlcPioqZ8lP5SVLtQK+e0eawKFUpWAyg
AkqxR2x6HRl8UBZkXcQA113P7dNuJgnmxkxS5tpTLZlTsxiy2wq1eywTUHuA2zyjmNKchZxGRfb1
K35FXnaSHwfl6ENNXZCY8l5y0oZ0aY0K+Ve5EWZn8L4NPVGWk7Yww4JbmEzoDgpWyf9t2iJ1QE/U
bJ6BmGuTid38nW9lQUTqYKnLVv/ZytzR9dTItcUKihcBjQROaSmOmvWbOHiijKk7NCkgIQMHKTGC
VRK3P4V/6pB7B/WA0CE4UqS53r5QAGc6k5K+BbA/Vla/JQibeHmTCRCULV1HnHF+KxKSJCAqKrEj
ZIYop+GfRpQhLCV/avanX2oorIT/QhasWXdUuKUZnhrej6RZupCE+Xf1jqe//aaKZu3nxUrUJ8mZ
5T62fnWSimx2MabokYLhSmjUYy0/k9dk204qTgNMeofdKG3xNDeo/KAwbqaQ/Hm6jCTQ/wKfEF/n
e3lOjBSBiLpB26mAJoTaU9mSAepZ5dKlo6FrkWW1nyeMo5tWpY2UefCyRwDruod2nHrM3K90+Ydo
TscGeAKUyvLKoF+v+aR5So4Fjf0YeFQUFYWxhKtchjuPEdatHBCIeXgF5uZnKFnoKW9oa493IkIX
FB1UwGImGwr3djEyQUkE0/esghlpswLb0ITZ1mzy0on/9yVgcy0TqZ2UkTo7l3X/C6TAlrF191zC
x4IPOABV+7fKF7b6YW0NlUFUCnKn6RNYpb1jE2jwt16NQZBhkPu8hnCWGsVmmu9BqcIUrxgw0qy1
RZuVcgTArGBYbQchB/9gLc4IjlkPWt4JvvgFyuwXvU6s23dTtNYGAWjDt8P4oMYToRvW1RNirV1t
x+f6UbiWL2U0eAvFNoRojKu0lirlv4SoASnIb33iER4vHZvoQ1P3mWGf5sk24QSb+lPym4Av+sVQ
6+w5h2BLkD1VurOvMGSohoA8iu4RNYZOihjzo5IxWzcqtoFC1kkwWBkKtJdlyDhDZo3JLdF4qJ1s
s0D1xlZlDv5YhdQaXFsX7OzA0ewrpvkvIIMu8eUXWshG/gFq4qwrpg3b1dynSzSpbrAtyK9cCheb
s+gwCrXJLtiEVgFv4C7mefC52xEvtyQOPzl9lLFAeKiu+kAUl16osLcn+MOjKuojKHeuFfU0ZDIk
0wmQnq/T05cxn47e1MdhuNgx6hu49wUd0W3MJAg/DyLhzS9PeEXO9cJkYot21EZAiq02Kz0i9dQj
KBDMj78ysZG64teQwYSAgQP8R2w+7nKPrGNQKvZ+MaFow51g7b7uSIBOWq4+ZZgAdi6fEHENkJYX
xB0h+M30R1cqxD0liegRRIJYmz3gJE38yLDoje07jLNTTQAUDdasXzeLM99kIqrT42kH6bDIWdno
i6hJWMX/adk+lvmcx8ReCDB09uKB/Zj8Ljsl6TAqJ39XnBvBIT5dKscrOJVOb7FJH7pRuL68o3Tn
oYh3yVcIKUWAubIVOefMjfT0OJ/QBcWhz98aPoMVCtJ9TVznYMpAjSKxSmEZHTGMlYgNm/OaL5Qk
kISa+kvlYSL/NalB+mC/J4tSHXHwdb2MHj6rgqxsBx3b6LCxX1fWR5Jn1ZTx2wNJ6IL0fmZ0Vdi+
v8YaazVy9q8LXj6pxYK+og2P9HjjTuj4KygJ3CtGhbFXdGhm98mRFD7WddS4sWjQ2cYabz6RxaNq
kfBbuWeiqU5ezbMOq5DS/3q02u2Ec2Zw7VnyZbRTxYuH3jSBDIgJ+/fb/EExZmwSKtx0jpcTy60S
bZtIyHoQ35zNkzVKxkcIB1Pgiu5VKselxUoYzSOqUcCL2UFrgVwKhJJpHB021PCfo/NvS2dOcGZk
dcZLto6+YIlDI9zxpOqGAhCj1YDQwNW3VErnkEiPjnDbm77REBzf+YPXcm/aqgBM7p9inBMeB6lH
+9H0J0NzLCIq6HGkvJ5pRrRbbStu6pNKQVJM+f/5cst+IOaD7NOvv42vSxF9YAE1nDCEIcSuhkJ3
hKVLZg/HR/TRctuUH0MIheQ5wgzGsENnUTEvYtga73Eg4ZLqF4elGlG9GYTJoCnmmi9w8COuLu1x
hVCtLbuzJxHv4WqsS123479Jcwh1/PilAlOlDllvx9gIBxgkHHQKSePnjNFcPI9TLrwIm8PzpzDF
UoQiTXSMmAb/LmaUTZJEZojTFfiEyi8O8AQHRvm7r1SYWAvh7kXa1FZ/2rbHdFNI351R7KT0e4nF
bV4RetxmvDamnX0hJCZ7h9z7fNPpfuBAjE84xKqgsAvlhc6iWvwB3oFbR8wqWV10IKqfjx66bsis
ts8GAo7bZd0PsNGZscsWshsAnmbGX828Xkpp/Lrtngos41F/tudHYvAaqPeFz4Tx1vssbmr41d+2
co4BxgWN5b8pnEglJKeuqCSZSzGqxjexMinljr4lhdL/dz7Yzl/P4yCYxHTOEin7VJzLgoZ48Mmk
uRUnwCa2qHgnucirL8+vA+zffu1DJ+IKKWVR/GoKXFJI0Xv4scJvszSY547AnXGeiiwrinentc60
ZUFAsa9L5Z+A2g0B0TT7izWmbAoTQGHgZ+QpxkuIMTyW9gOn2Com6jTGzv/uhKG2XCZWutGZNWmC
2m0q2UYBU22xQ+GRSzL1WyDBgVUMxzhUyCI0uUhRSUl0X+G2h6YOJUKOwkp429AaULyyFYLxZJpo
DaS1x1raeldmXF3ROkmkXBNf6//dcU9oy/rR884C93w5xVpK8d2Ea0wb/tsuKO4tMXdvZkWNVa9k
bK3hnq5dhcUWFTUTEN/PFHGjK/oMtLIKo8rUBYva4iJjlQVapf4hQR6eNj0FgDszdI37661IPT2Y
SjQL0b6qXSPtzr2wlyvUTMQD68wdWGDPP07lCTzgHE8kUFE0N+BqE053k60Hio8aM7CzzYcXNZbu
GcqI6toJDuFoOZ0kpfIWymoiSv7w8XhSkHpLIRThoak1x/fo9nlzN/H/0pUF/o1ed1U1jJ+Fsgx0
WukZeBAT8XJcgPuXmPK5sRK+7cttSOLex7xjvmiamPYvNBFRNATWxaiQUJmHI9hiWJw2f/E9kJ5f
ecGs9+fRnJr8uUsLfdZwJZ5xXmNvwks+Cbj+GQeszIiWkzotmaOzq/goPyzmVwRYQTP5M9+DjUgl
8pkwtyoSGQtrBiykNfXGwwOn0S6xRSmtsHF/YA0ixmh2aq5IR02A2jvXq9+Yf+4yO+qhdKRqAkau
IRnFBL4hg7NZRnyZjYqXLp0mUVpkO61CJ2tdPc/TrWXFIVyYqPU4qHe3N6FOcXQKULaRfI+QorOC
tQ3g7e1u7zqIdQh9WxQtK1YnNim+6smBh68XVFv51oG4aRYHBwl6x7sXKvvBPIquk1QESEkkBVjg
Pxc7sGB83bVl2LGBNSG3f6bACptiFYrT9CMFLlgpTQBO3qUTMjU3Cj+li+WZYEno542KZepLNY4K
TH+p86m5ZqMmvWxMXUoPMRgbQNVE47Ta+HfePJgZyUnqQh+h+4oNztkIzIykqmyknh1VcrMuiRsL
Bb0tzyvOyHAkEm3nyuxnhwyZfmGIviVqeUISr6CngTMOQWDJSBm0MKLV6X9XkQrgGk08mPtro4Aa
2B2USfr9vCFbDbzZzeAr2Uih09xBFk0Ze6zptr+jrzeqTBcXbev2e9TPv8evo6TSapcWm7JX15w+
EEH35gMP3cVzZLnY5c1V5b1loaCXm991Jpu+oFhu4PbZyKXlliGqaAMI/jyXnRQmsc8sKrBmc56r
fMuybse79nd76t6wIzp/xiWZ6L1TnMpei+HQnYJkkxBOVR8s8V4U4WF1sKB02sIyFjf0QgfJvqUf
AH/oo1eOQg7rFyaxMpjaBOTvPX2pZSmrGq0UNrNAvUhGjIdw5wtdSYFcjV++7XQ/8KCNTYjgL2pF
zNcawE1okclosgM/iO8PV4p5QN5sEfsmmrvqXz+1VXFtqQkOoYJ65C9QbmJGcJ+JLj/SlP67cpWX
YrUJXYTvAMQ9d0p/mRl/92Ld+OrF4QUJSCkWxag4ddDiwqhNGDnYkGELksXcEFjIlmge/dGvKZN8
kX+1gVKhlNONPNV2B6SvotfNAFinTgfEXRX1fv6FgR9b2OWUrbyezKID/3JrKmqz0OM3pMpOpyDY
hKLKRawbv6D8/tvTaiKNnrRm7I//ImOV7XTYYSouhfuWfjSOBwy0QxT21+O+xAs1kggrkyQfoA47
t7zgD2vmj3k4XxRtAOeBUNEky0a6FLwn+9hFP/jQCPLeRVxgsgsgJRwfNOOps4iiWR8gQjbjNby8
mDieXNMefXC5S/q/3ZqkHKyfz6MYtoviXTSMOIzTFIksHm0mC7p/hmQ61XzIlZzz5dZr1iIjKf4I
GqMirkRWpRmk4DStW9hjZtKJyAKMym2lBvDI16mJMOjaVermfWNg6sShz3tp1/uWO2PEP4QLblD7
ZgQjg2ZxlsPdkhMqnoJtbmO94hwY7QQ2gSDywMLx4rvvGK4jUboPOrQkPgL0QXp8YUXMSEo5Rexb
IRgJ5n95fJwx59HAJzzgBmpiOwQIZuE8bZmYuSWsbMDJhjFEBHSS+KgV1bLOmXmpZizY8TnO9avA
/VfIx+kCWBvyEeFvZb0BhZlkpYW8M19LF0/+5I2C7/PrwQHZCeO49EvMNcNS0+v5O5wTaopoqDd9
EiSjFk9psJg86WYvZthwkMbffQ5KQYf03v9tdr4dz6luf8pSkSAqk4GK1itjrdGNXfYLh9zI77q5
3LoyDiMC0ReaTroO/zyh1n6ibkTxQLLqalMjVvmEUGASxnUi1BtOyObOid/kZuJ2CD4g9dt7OGlJ
iDGHQJDwmN64FSbtEowoDffUO/Fk6xnHegaE4Fl3cSW00esqnfFFxKmFZR1FBzigmx4LmDHFP0y0
P6N5/MxlbRwJFxjKyjf6/L17iHTFVKUrj+4KjpUiXpXQzd/RhYSpRFxPRl1D5dlpaVxK7533lLWi
+cXMfBPihrGV79v3OQByEcKI0/HKwofYzsU3ThcH5ZZYk65gQF10IPCk2XuwdtiaKzigvfrSSpqQ
0RHmdBhFhO1MhKC8Spx7dJDclMlUklq2DEC1V0uTvuaVPazFP7kOnxiJAvRWcAKqqHnkh4mBorcM
bbgMgpIf87loaVXu41lqQmGkHBhh6btXjE9hawOVrDCD8hR+S+mRTb26uo6TNEN0SHHUbNHqoexc
7SYfqcDzvLXIP+jQr0cWlFyLnCBJ2/4UvHafifEcrn3s38MIR3Sh+yx9CM4cAUokEGefDmXilLpP
Bg5LxW2fllg06el1iZoyOf0xCWXzn+yNB5VdJaVneNtcYTwa3PZnB/qXunKGHokbaVqY9fTp5QCO
9snerUOJ8NJNeYfoK27jxoBcKGEkYpaxLvujAA9PVl7PX0u9G+bYwKxbj75/Dv9PPvwm66u9dr9k
+P7A/xbYjMkDkXIla+COUSaQWHwn6M1HT2cOI/U9rCDDqch4QNd03RqMwXmJMtzX+J628Sn6vNZ1
RUnPdW5kODOoAOfLutO39VndiMu0yb1zcnlFpa3x1P5pNZQyd1jUPoULzZz10BOsBD7Ya2vahV8p
WzMd4VrJ82sjhjQsoQGhZa8ooPpRA/V2ihDj7f0yVcGuPYYB5ZyR4Ifet5ilHEjtFAbkqrzaYMpC
sFMYKqM/o9Vv63N/XLlSg6gzzUY8ZzdTOZ8IWq3n6ShnF3xK0/l2ccU/hRz8ksIWTMcvkBIC6SmB
bVnxQ5CVFrQOHmoc79f8sZTRVibiwEJUhGRxcaBbVd0IGcjRzzoXRIAe++6ZlkzaSSNd+OW8xt1O
DvYQze8HM3195Puk8cIEhQ61/yebu/vMUn4vJLCnkE5pJhwyfj6EP27U4oV1il0atQmdbXHEyC/S
EAR96f/liWmorJcB5plJxGxbXTG312Adnvt5N8MJxb4ilz1O5U5VvdEtbpQbFtiaEZDX+fsbS6WV
eOM7dGeocVCEeS7Y4GhQMtZphqFtmljxSO5Yfqp82Ani0e/7D40nmLjmnrPRmFlpFZ74zokvOu14
szrJBkz1u8+2fR4VlzCsUCpaVx7GMQ74BS56utzmHNrvEaBH+P/oxTrbOKR3jd47t+ZK4/0wVw29
qoHE/53G9GyDAwHivEdPqNKSZ9LbJzG8oXb+bORpMgioAvVIvWusUMrDOScRr9iq64SfomU3ffD5
Yi0MQgNMgC9Vpu1ASDQ+Cv1cRaoaUw9N3z70zytJEWg/PPIDmuoIW381uqVvQnnLbfzTgXmeSpz5
TabQJJw4O28kWHGJNyygPMCcVapc8WX/Ld4b5NgnqXwccfwuP18j+sxiFLyd1Tb2qea2+cMOobVf
RCWus2sNeVYUSjuS65XmEz80H9tVodc7v6G5GZeGKjhsdOiE+NSz/7Gi62IeGfZoXxRVQK8h/HIf
cQt5v55o7U7HKCtloJnyceVuV2z1m7iaejI5fJbF45uHj1GdoXUD0t3pjg7uJ+sZeqRfY8AMxkCt
d4uC8SFMN9xhp12IOayefi0FpX2QsPDuD4xDvDH2j7UkNBedbimrFdIiO2crISgxA6SyHqb0ViwM
LEyqFY0FrXimgg5bDIsKyOmhJreATl/+vSmUiRiBQx+fltUB5ESpSci6DDRKn2nq0eyFtGMlDUHy
IJwD+ve8UQYcu/hC7XQ5xP72klF7xSEGAUD59UfRc8QRPKLaoI/yseZNNyYdIPnugt7g3o96fN7c
yNJrlfjjHLsbGjGHmhPQiNFsH6i/BJ4JbbRfO6usOCfoXzoBnb6VU6L0vEFr+ksi9lhz7EU55P0g
gw9mBorEFuBWaxYLYV8hkfJINnObLb3iRmFS4c05AEMn47sB1hcJ9gnvYWiLdV9KXnP5Dcww0lhw
tahs/b41DX4UgAx1xTkzE+68FD9vOGoK89BVN4uBdF6GK6GMbaZaX8JUxOz6tAPgPq3Biuk+vGeA
oFYXY9CS3FhHJqvxR6OrEv98GTy7+/pPX4hL9zjo+g/1gofDFsmQySaQNSpN3UgusX3c5kasyvCM
mKZJV3teD2Fr5XK5HqZPZzuO8otiSyBk7cNXCmqZv4kQbXw63FfW4E6ikqcchvcu/wSQBmza3WC5
7H1cbcO3qKu17GYM+a3yi/pdfXVGOmjZHRh3NK3fBtTfc0FO9FTIgX+dCL3nk4mvnQQX9RC2pe+B
4BsuhP+J3g1IuMT798ignRP51+Q+BXZ/CnGlxDsUNc0HVdL7Qc/uwUZPcVozoFdK+ySfu2ZQe9XV
3vMuyzyazMtp54t4SEHGGsIC6hRxGxOqJkUdHrB9vm9jIy4wrYVd3smOE0Hkqr+q3Vs5WlByfWut
cXHIZ6D4k25HhXPC1HYPkn4hOSbN8/IjXVbnKU9R4Ffa4imD7iBtcUsCIC/ro3g5e6QZpzM5fJBC
u5d0zJX4uINjKdmaIhfPOPc/lE0dNTtjjiyEORlqSNjRcMDljj6+oPOeOc5httNo4Q55PMLiKBAo
BzJ6xWKhTDPlZI9P9bo7Qa4ivIb64uG5Dfw0KUfDtgpcqElqUxRCFnePUfAzaQotgvdNilH47bot
zICk9AGiV2E5TJmpyQ5/avqa6CcRV06uvB9SgSxnvv4RzC0l4eiXNIjo7VOogUhh4Iiww+bgxc+h
sY4nHqrJj+fDrlxaOGg8ADpuHmw4Xs5Q9LqRqN1kIrrWpCpLI69vB0/hJ92PSo3qgIlwR+sH6jFw
fsON0eK5IT3TMBzhU8MhVNSP8o35/BgNnzW6jVXkZQ2NBfg/bM1+AH4MNZ+gFAEHjR5qIJX5NpDn
l9sgjeYfuRob9dkoid8LqYcodJfw+TbHUrMUJQiFBNr42EsWYipMXbkUEjXzWLCerY1Ksm6VYvkP
FsskSv5GPEOwg68eOVpiUUSBy22ANojqo1aGojxSSKOvSAhb19TKyTRhveYT09wmN0oPBTqu2TCN
ai18/KBSHONwWp4QDF0vMWgqTCfbX+y9K5NmF3cmUVZLWKFw4LN+ADa6YqM3UqA1M2nm5YdT4vzM
6bZgB5k22cJngcqm6XY8ZRKUJ92dqXV4Rkr8AuGisi3LESV7c1LkisSp/m/WGjYJaFNhRwPRHPye
7omTVSUXkZL+KdoIwdSUSYopZnUK4fcy3K9tmXLrSQFVBlQEYVxl8IujFeXFL/5IOP+kCrQnRtmD
zZH30eU3xKabBoPKWLEsju+tBbxt5li57V+AypmdscNT0SLkkmlFtWatmw00ahUolh5WpG7yHITn
kovlvpf+DGEOLXvQOzPz11oZ4TigC1YI4tLHWIaLxYg+Cr+gcjHsH4uKDoOGJpzBZ8/cK+S1vK7b
EGY5Ba/+gFamwrzIga0uvEfX3elJDLbo1rRaOzSS64DqsD7gbcrI5476CCrLQJcuxsCcta1rv8Mp
nkBkWrfcXjaf4QnSElpxLbKHblbaqbYBCxMv2jz/zYTaXp5PYJfeT1a2Fp96SJH5ShbKD7vUh0rM
+OrVlJUz3Wb+gtGkN1OQQZ4XXx6GfRchmA2i75IzpYQBr/6F6ZZ4+muFPTn5V0ql/OouToEdvZ2D
ibmVlvCPF9QyJ7FsT4zAUIubsGmFKRxYH+KUai5o0KJ/JEwFTgwbbaPJND9UQnLqGpSlRIyjgJuw
JWO+VOkYlaPbA97JIq+D5aBDfzSG9D5+u8q+SHWMoXvCZxP+x4zVAezikhbBPGCGkDd3EXhqbvJm
JRiZpNYi4RaNWVKYrlo8S/sIhVPuWzf3+HkygD6N3wb7XZrgR2uNA4KFS3K74pI/84IKibWtJHr5
jvH/Ic0kBK3BjoIJk6tkyxXsCQcrFO06miNkTLaGf14PNMCMDj/4UOd6w/xT4bKVXVYqT57/HBmT
E60HocNqAHyOgxxq//qw/SZiplbuzEDlzeW51+bMyxBEVM2hOqld4403wxoUstvDZSqzQfuvf44d
Nfimq8onkF/bW9a7qhyyy/Esr9vRF7sBzR87ErawU/UfxUEp710Dzk1h4YjItJirJS8VI2QtzWtQ
zHODVB6kyYYhlnKen5NnLSsKZAMMXEUDZR4dgJL3ORE5QPsmzZ8r+7n9LVlmRIElWgEhi2tFAkXb
z97B+2s59WwLfWBHcUgLIJeCdbyCov8eCJ6ZZ7m1BDkc1GhUtMl6nDikKgmxR+gdgW+BodhuhD1O
WkNKpOOmkjxeHEqXQ8YQPXY8xWbHL9AnpaC36A4UM5OKy0sliL87LC3QaWyEQvmjXxxY+ndJwRNh
56UAbQW2fqUp2FE226tE063WORJZfagrIYJYEcPFLXi83Z7LanmWKS6prGtxBfHfJ2rt1oeENpQu
GXJivLir0PhZMH9d/rzVx0NZAnHEWZwK4P76LV9v+cF+g3c1bpJscvX1StAiYLsjv/EV4o0+Y7YK
bi6NZVqS08imrXT7sGBniTAxO4+sSqGfYiuiUsS4smyQGonmZn/JGeqDMLOolTVQxWBBuirbNwvm
MrehBsMupi4oDvCvY7xd48pkQhK0YfCHVI0ASfbM8YLPXCYtXnB1ZQ7r2CNTmlNoZXHIEGs8Hynq
LXSY0MBXmACH5aJ8Bb5G6TYOGA4caVY9BpFJjnmvPYPhu3wFIfRqT0ghOs7GGWZhIqUdFcST+vhY
XziiyHQF/O/Ftu8HiEvADB/i/cvFM66hv1wqBj6LB64JaX28fCPMk9lTyHUJBCWCS31gCuE3nHTm
QXsRvkZWlXQe+3YwS1YBUx+ZZcW/rQG/I8evWq4S026WXcDnZgza/Bn6SS3VfUGbygG2emE9/eCw
ivtHIvbTuRQzcfcXar7FAkeEYCdgCPbwaOOUQuwEkGOEhBrBY3yZHGmQX3D0/JnOriWpbub9u3cp
9RcA0XFrgQoInpuSxM4fWRDOk7rXBl0Z67j8ie3kc89yfrTVe3uGTGU1Xx9vXaAfvJUU7Le7pZmh
pIlw9R69kWa0XerqVnTb37xmZ+wLoeEMHlWmLe6wh02eQn93CAgCds4Pw7ecJMQQUpYC6ozq67kT
ugUvt3Cn9igH7Kr2aEk73egIhjwimhIGBa51cJWgwUyoOzJ77ES2yT40EojO2YLHe5vHIonDSa+3
Ir8pM8ZusrE3t+8A/anenDezkDfB8yUfomUs+tHVzSpssjpTwl0+UWlLLGmPlf24czRVz94ggGy2
8b/Bh+0TUMisG3u4ITdkrr5cE1sAewh5QMdxAfiI1YmGbVbtiEpIEODf22b8QnaL5XFaYFPs0mKY
zD6U6xybkxb4nMW2rvSgzWInkdCYU8u4ApXQODLHA4IYJCGFtl6n9ftw7GbEocn5D6vE0qkVbK/r
51CT0LzuNRK0Rh+4BCgm3HnE+7PgZ7NxMWp4wK2R+Mv7upAIgG02UPfydlQSGIjNFPymAOJI3Xgg
Lh7bFShaRgal3uKxyZKmp1RM3X2d7F9hf2JRcIuZIsLjrU8BuMcEBn/4pHY/RhPoIFUWL3sBJEZV
qKNZHCpjBPOB4C549y+E2GEtHDTMfjx9wchiJ34lsOJE2KE4Hx+1Y6VGw7MqDMpDfnGrG7q4PCbg
PDHPhgYYf2Uzt5jhRMrZKRUzxXU1LwRxaMvulSePL4ZP/CAxlVqnVGQKderrDb/5ADzJuBR1MEZ0
aFI9vKnDHggdpvD90q2rPhYEVi2k2CfMN4VYjUsQo9w7ZCQnNcaGsbXV5/EE6yofSruqSmImJKOV
/8DVJ4GcflYM+liavzs2OGFdFJfuBbiKoDWoM1uXiD05HhcjQHuFqVuOAsc3RBrKgf1CgiGUIM0O
fjskl+358fAaaAbgOw7fsWq7dKMYhaXLrZ7iENvSbkpM2h/PpONOtPpeXrJXbVGBifBZj7msvLbE
54wMX71GLLKlwAnHOV2Apu2+OecKYNOEon17LN6j/i3hxl4+A5XdrTX0TCbZk0CE58rbs9MWOQHL
qIeQrW7FLxZ0gmEzJW37mAZo74YKEKZ3wNESd3s1kqwFC6v3NeKWJLJwo2VSfQAdvJg2dRq3001u
kcYhQYJMrMTbLl/B9R1BHfUPalDCUZXr8PtX79/j9RKJ8I6AT+ySOrSbl8l3zjmNHHBIGaVFswje
CcxwtoG5/SDAtygLkQMfhBAWueznlmDHEAh2lI/pb5CpngbVFeDg8V9WWM8OO3q0N8QeQu0JCK4N
4a0ExUmZa1Uk9+Udq80F3CKZvm0A6gObAfnnX8TknVQfLqnQtmNHd6qm9MJDA7TCmOjZr8Q8Q/eo
MI8WrdqDiy7OUAzesEG+do9/ZsHC/kiKXjNLyLILEQ0usTU7Ip0x2wnaAVmRcu+2ShdShSiVjYkA
a+VYjkSfw728rnPVxbO1brthIzAY+iaWl4IQZfUWu/ZUpTKnGN+lsA7XSxisGTPXYcNZdffDGoK0
qdN8o9ZwEkgyfaNbMxjt9ARhuqJ2SVL1215yXCSvcRqz+xQp2O2zWcC8mcO7h3gdKdGOOl+8kQJa
x5PnCAYG3KaXAmC9eqVSKguam9r9h438Mrv/mnPhhlGrXcB0XBfpEW8tSG3PvhPfCiakec2CuII4
Kg2g4hiVSzOCHgJcPJupuY8HG5mGg1f226Up8EsMMj9lx1tsCLqZmcdPftTqi/Ep0a+5OYXnhQ8r
Ojjb93AzSSwSN57+K1T+txuwNgFInGlhfiyu1ZKHlE0RwqoP197meDASrTX0DNGCwEs+/o7T8ngL
xg6BYfWrG+Lc6BcQs78pM9AxVeGbmABNdm/xD0sF5zqNCUmnjrutIel79SxgP6mIeHklwra/q5Fh
Eew1j8NnHNLFnfAYsSqIFKpfScZjx3MvzSnKd9ecd6U1vubJAhqB0aPSeC2KT++5JvJE5JBUVG5r
ILNboJrTqL9Nsh9mUm7FTWgdMi6QybuXbRIVaIH0kgOGiidXuDMmOhGu6RZt/tJX52eqjch2vDJr
4e3It6GwyOgCJIFEPUtq6Of/9+G/SsRzF9UWp/DwvoHs6lqZyHoQmSubnAZ03qN2iWa7+WmcjDTN
pXyNbKC4rLfB7fa5TLqcxc2VIh+OSusd1g2kxlcMXS2R2SRnbtt3PtFuExMz/e9VACzpbWR9ihA5
Liuzlu8EofPOdmEfKpt9bD98XlNsP52/5gsIe0vLxcSvUDz+b5/+JRw8jvto5NOrYzepm6foNSvF
jmwFnLS69oA39ZO4ibl36CJlUaNvQfxWvFBIQ8kfcvXzaqg6g5rBSrN5VdorpdN5Te/UZr3/qgOh
rH1EvUP2gCkn64Zvg71pXctGqRxiHbTQtY/rQ3yvq0mav8W9t1IJ84Ry66z15GKB964V6Xd+yK+H
EWP4fJwfhTh7A0QGFJhT60EpFeAlMzPnZlpok65YJYWtAUN/4ULJ+IfWdBsmE6YZUgqFoiOWWpsO
N9a952l1S954RK+hrV9c//h0rrzZs0qdGFBqSlXD4JQSJCcM5hBLWfXCX8zJbMWZu1Z0nYJyXr/7
wfUTkjL9lxs5t4Qgd1mgW0hXTYrsAzw146LECf+oCHrbc9j32BVYQ6LmjQYTc62I5WL/EuOn2zxY
P0cyfXvse7P8BTNQD530p/CCAfTRhMFC7eZLEjQ6tBs/Wrl7k+AFCoT1932tG52Jx23sDs4IH1lB
27ok26GeGrElgWBRCRRuetNxzhHUpLfRdl5qVPdj3ilJ+Vy3Vb1GRj0+XeIkvP7NS9YPmSutjO6k
WDqDAGJEwbsmuIeHBtM2blKfNMd6H0fYn/f5hnKSID7vceO5go3WHjnnpG1jnCnojq5OBxEhXhPu
OxATjzDVkWjAf8MSrOBvTYevyOBU0U4NoDoG2KS9xxn4vSnKkEt1FkD54Fla7N7Mzz0J4NGdIJ1J
8A4P1YZCshzT2dAfet+QKxj1vBBYkprxWsaw8etenjOVzAUP3MrZoDtiv1UwArGTSPLbFUVwMU04
YlsmHXfxR1u7gW6o0D2u1zUGNfINBHWy0Dc3hGvNfY93SgFEwRfVFuNiHShh7krIHNBb7M9mGaY9
TtEZ19va5e1N8Q/+APIWQj+zVTNgkb42MO6xP1IXSgoogKycXXt166paGspxyNXCo2W89U4YucHP
QbIxCwNPcNYfU+ShixbC3+1tZXoPzHoez3860m6aUE0xWzsMryhYJ3POnpNHA9ln++wte1K9onye
aJp5KaSXhdlBH111n6hmdjGczW6G3RWv702pLIpd6w3cMRedY7Tho0d5vzZVdqqIUB/pn5UvDYtY
45I/UWeW+Zq6VEpQZb45vJ30L1pxvorm9rpcW99hsl65VuQ8DEjCTPNIClXGpL18q121ipVTPPBa
5acY/yP0S5wTkfkW8ABBGWdlHQHKRnAmn5Re8W3dckT4k1P5dqxBeNhfTm8MMby6sjthirUVS9xU
Gmly5/v/AUjBGbL5bm5qpd5rLDbldN09+mIcPx2MRFNUCTnvg2ST2sHFTTmUkzyzoW455x9d4xqb
MztMl51cd/creVwijLT9fSufm6anmL2T/JsuSSSxNckCeA6f87PnAM2Msb1a5vIIUyFYTQ9f0+bn
6BrRIHflw6lN+orIGvDYSio11L9ZB+DihDfSXIITIYEiTSOHkywWpfz+gSyJc7LmuxzpCRSAMLCa
rzfvdnlov8eQtcyU48Z9WkuMj/X4kXXBrDTTRD+unjAojo1LhJBc89LsgLnX72JBkhy1hVUwt/uQ
Pq+L3dMOQkC453/SOREkuNuowApNaijgHyYETLK98yn2myM1SIdozXaTo5C+8gAYnkge78sqRA88
Z8zXy0micviV6G9So0vAi3fO2PK6SY5WGG41yfweBij9UUSJ06DEf5e3esA87TJx9rtqaJ4Hrtrj
0D430devdvItjknOTSPHQnl/gE47Jf35aZ9MVLvSVvUTA1ir9VKzrIbLgBTJLwsYsObXo9XA9QAe
5/SD7+aEK4aCwDeUsWHKVoo2mjykN+vLsipZEDqLS9PgmeHyzX7Bw+uZZ7GNJZsBZdVTpZjMQchi
oB1NVQ8jRNPbpxaPrTUI3u1zj6HNEs4r4hc75yMDCywhVBLa/iBG+/G9JqdbmHxO6jT4tRabvPg/
+VjQFWYz5GWDNCf3R/uS
`pragma protect end_protected
