// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lduZDlBsPMFVJrhJeDstDg9LfNWNUXj1BsfgC4+AvaBsnC94SmGT+rQhFgSccmF73/B2Rpi+LWqA
kfDoRUS+d64DBWPrgRe07kR1YV5vwqfrJ4/HViGIHT+yznbtVsmZndkKyZbWQhMCd6IgCxSK/L86
Z32znYdWAfGALhb/h8TOY6ujBxRYE225U0De8N2ni2OPAvLeIyTY62UpffXiy5I5UQtAF353kt9P
Ly/lJQ/Q4u/KbnyA/kxOYb60ZCGrBRAFHMJR2c/LFSVA/gYkcWSQPwWfp83jY1fDr0qnm0oXCrje
LJKf2Ra5iJwVpPEpBI3zuSAVRxNpCD7W31iBMQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Mw3gwbmktUnTUn4MRWnPnG8hoI6NW8S6znNjvnIlrMvHEdgFMB7ST6iFcbwvp5OoCHb8/6sEqqcG
mYy4JdKJwyzHtJ6T/OZoLVID+4NeqCZMvIwxu7PPu9kLnzUjQmJomvKarEMvE6rC2cnTXSF1AVoJ
BF0hfkpNjbz4tB1wFOs6ZA/fglO6CpRhjsGd0P1vGszABYh2RhMKy5j+PlPrrddsfEwV9kJTyvRc
t6PF4qYzT94lAJW65RZTOLT8MTWRDGoRRi7yxFnbnB+qMhNlTvHy2NqAOO0KfNbVJznNyk58W8fk
06iT4fakvHVF2oMiJIX9/66bXn5pdu+KLy+KTJNzO8HO0wAtQNVOVB/nPybVW20IdLbNkEuS8Tf9
auMlJz3pzqmZ3v5RfkJyYdSvMj11JZtNNtbjtS0hDFZC/ejmL7bi579cHKA4Xfk6yrZ1g6t45/iO
v2CjjWD8yeeuz54fW7zhgt6K7ShYolJbZaxta0ctPryJkLV6GDn8M81/y9KwZ5q22CRtomZ2Z2uy
72JGyTAhEPJGNa+ReSr6wj5On8/dUFtQVIIydkzNkRQMjvI3bkMlWaZUVhx5Ojs3BgOTN3y1cswS
ZkzYHxjI+Xnte5VhB6r1XB8QXkip3ClHqI0nwXCd85cj+LLAu7d+JH3bInNhMFj+UojPqFhvPBUG
zrnTMQQbjeI0Z4WyBse2675GHm2VfL9Nb6UVPvQK33xKKiWFVDqhmFOOHMA6iOWW04GEMmOgS7LQ
KllLngRAMhEeZx/JK2+Pqf1OV/2DFY5foAXNt203i3CFwRiW00gfpEZE5XVDbIUXkRaI+JVAF3yy
LEouDG88B5mwwwMpzC9lO9HX6C7jKz5rqeSaEx7RQHHeUDFN0gFRawvdz/NkZcA8dqVfKLb+peN4
Wq1dXWLn01noYgco7ayp+lIV+nvEVyY5eurpKT9RhCQ0C3EqRPheMLPyzjenkIGLP/AqKaJfOi68
kcYSUnIGgRE0a9PB3SwCGpSe0oOKA+hr8RBfcvkvPwRUvefhwym0qg/F4l1/Dl20Sqpa9NfPM44/
wN2sH5ucqmTMCSZobmZpQRInA2HeSguH7SX8oUvTntQOqtjYUVkHfxFj+R01FeuhXAKax9BlxLX9
+EKcZx+ThERcw+0XoVD2hbqHG6ZyeV3txQmeFBkkUDgKufKdMQ9X/n4knapSdD3eP6lK1uFXHZjW
ajZlFTveYpASmDzWdruXJ4B6ysmuzB38IJC0mPT2pvdHwgBq3QT7MKv/6uWSWBjff2hjf4qt1dDj
S3SkeN82zRhb34rbDlx8tbLP4+KRf7LWatAJsG2cXUsXeD96hTPfHM9Yy9foWIJotsUg0DLsZ+4W
qrTfNuI5EbXZmrkBYa9XI0RNE/o9WgLNix2NJxCvFfW7W6BHMpum0cJFGbbNFr23sX1O/CAkr8Zo
lBRz9l+YtIGF7KlXMmp0G6DGpItcPkyErK0H0OHpJ2taOsBcCLjG1J1/7Hrs3eSd7wmXAJbVAiYO
9dDvhja1Wu9ViTQ6Apt+Z2Qu6+2IYkqKRcS0pyl4A15b3ao5beEx+sCm6thI7HNOuwHrgSz/c+su
f0Ec9GhmP8/xpgWHL0F1MtX+2y5jSm3rxsVthGH8RYxn8cwJ7w9m5nrCxycl0tlYpA3xf8tpvtTb
Hj+xBLvTmDuuwI4I8VHzNoH1GY6eRrTNXkri3wrzb+5kLCqTfcB9CRH26alAgb4fbf0PR2ca6Ftm
is0W9IXi8zgMUXGhOz5JIuYf5/92k/OKNLf8IBoAlvFs3Cjl/qNUt8nBy+FF59vfxtHo7W7nZAdX
CuTEUUmYlmiako82TWgq4bx1ivOSSkHGHQl9JcN06tRr0NeBDGuI+IP2QPV22If7FGvmw/ygeiZj
juCtKQmIy0FCr+MINcOHJyCIMv6/vFpkoLUYqUqpJgzPg9JZLK2BQvXvz+ZUOSr63mg7kJnraIak
CjYRXIutYWo3lHMKsLEzsiUZZsL6V2WaThOnXWJtPxR95PilIytTjI+xWCliRWY8wdEufBwHb9o5
oqjJCPpE8wS8PTh2Dylyipy+ZZLO/ojTwdRwGpCbyF/8eodEul/1t4g30eANQB+nKxs+FSJennSI
3kTtHgDU82mJTSXahXsDBEhgAVUYDKyp6yK+aCw1AC4Rc7xPkimWd7Fk3wOA4GkrrCvBzF5pBaie
aQHUs9exiQuDaZUqBY8EOwMGsFROPlVF6v5lZC52K+B9YTqzreJsJtr7lmdJYAX2gNfnGtogapIS
giSeX4vuLNEEZUK7fYhJpzfDBlTVKOfKsR88qJbvNDO5BZsISPpIXp44FtIXQCTNwhLZMqrBKnHo
GW3a67JpHd+cFK1S3ymE1O1k8A9U8sg62BGtfMR3MLTEBjvieydFsQMcwIOEO4kSrDIz5cESYJk6
kNX7u4wYXjlCgOq4A/GSbIEOlR9ZMcVufy93rVYWaicAC4E+zFzNe+jCgJM4b11RexaTcQc1zukx
VtAOHhLGESOwnZKxwG93rppo5AslaiH1H8UL38l4ZikcqbPvo075GlLEYmTtwIyXbWOSPFUhANV1
MFpg2DYQ1ujZGKlnyUK6eraCWXVX+fVbylhq4UTm9eq7EGnRj2uSGhn32xa+4gzXR5gJfbuxqrQ5
dFDXJhEPDNmkxWrlmUCoZhyJ5ItZDwhAsFJHQ/7NDSHRCUrL+PQkJMNd/9ttZi00/50y/mlXNUFM
McBYDYWZoaOJNjkgs0YHyZ6+iEg427jdiFJK79OwFQhhY/AW5nmRnwf9mPqP2RkmqDfFWfgd4QPc
AHGYastdtzf/M8TshZAB2mSpeuB5nVRXUNra0Dk4Xj3F0ZgqyeSc0KhmRRPV3SMlfmk2Q4qAtHZA
zeayhOOo4+wkZCdx0WbzIlp7l/vvVc/idr25zFRNrgYYBoPoihnIT6wk+shmGrMbUfhmB952TN43
uqz2SjDKIjNTiIlHbarUohqW1jwdWCNH91b3zMiaWzo0ltHYPC2eO8l5IcyOUPzRN0w8gTVPqCun
uGnQ/zBH/huDWzrN2iKpjBdLix/DRkxSNbgtyogURhPCRjEaqn5I4UurlxQAhsJuuiw1jugHZDSN
EDPP373Hw8M9DOmfHomUDVOwk0muSi0YlKmZv0ON00P9CkKcIM8HCNzhhaUgr/Wm1ivCzdEmcFr0
nSZIylpXXiPCJ0/vfnl+/5jeiAaRZS9lTLQca13oBbpG5SFAV58qhMP5oA6Ke33SbYn54PLl8UOj
KuKjjm9Sq6oWHvlCGtyjDXx3Xgx1jGsv5RT8S4CWnVCdrC4NjUxfwOq3d53YYT+S09JxrSWkDtLj
Lfp/62jcI+nmzQoWjR5cIIDLS8PmAey6XgOumFDdmq0eChtaong7uU/nuW+Qg7Zywv2SmUYBpaA1
O+ouaBgmRPsuXBHvi8Oz3l7Xkz26fy4PUE8RIBOGtnsWNLcxoQ6dpoBoLHNME8xKZYmlV364svgx
N/eOAvhOxbPJ5/c58DjnbrmukycKoDa6IL1lrl1MQul3m9PREdmsEUuuoluYpfl/ddXBArdlFDHJ
Skpi4LIUdwIQEvNhcjJgeesK6ljDm8WJ3Irc1h3pYyqLH9QjIemPZef0TDBmzXY/EzZbIXmZxt8z
fwottJnpA4cc1yvdW22c6LlJ/nTpbi0HJFBrjUcMGch5qYpuLufVddSB+Wx0e0PCDDs+22UJCQvM
YVlu7V4oXKSv0QUj8xK9wYVOg9WYAj5FFv437hEI2zdOIHEneyd+wpN5lXri9GLrYGX+zWdzdXwz
O0NSlQ/kkI6g9O16IgE1OaoMI0t++4mqhp+Kt1Nz/Y/v3YmF9yFLIfxPORawxobo0g7XRlDfxcP/
X/50YEwvL6QwqKszClLVTNsHSrk6kqCP80tU/jRJ6tmnzsFWiikiDtG96YVfFCHIgg6e68cN003q
Mit2x+icRz6bS+IvF65uGZPHjNke7zXs9sfPTUnD04NhTzgPSeGlXN06HDEit0+TEdsnkStTocBu
exZy3rLY4h6OLBib+pkPcGq1+UuKKx9jL3Qw61oLEa8zYYkLoX3u9IYEp+vMtiJGP9xacyN4WceB
QJj2E15TkeKBqx3CF6/rPX4hrq/8PMXCFnm3zfB4g5rOcb0jQDd6sfM05gt3uB04ZISLBydFqw/J
m+IGs4GrgMmA5PVbUXALCwtXqg7vPOz8WI98dbehSijTZTDYAGlN9/ntRWwf0IHtRSJIlHxxwwef
fWwon2sAQsG7XLhCMXX0iaIPw5DRg/HUo6/XxfQREsSejezi5zNO8dblXc4rrVL+QBRb3WkQu1fQ
sj0pzJng0cwag3adfHf4ZEsnbtrVgdIv/OaEE3uQqR8PLx46D66aJ2Rf86078QXxVxCswEjyDCHG
yV/CI9mjGBbj55UqKcM5f2WO9Qs1BW5GcDByPeCGMsYMqaEVuQHvxrOksOOjoJ20PtU9Qd9KYlT6
7TIyi6I6IOnyOLMYWqS7RHjvLQf2oV5F55LYMvIbydvFJFy59d2Zcu6YRpTTEDM6Kkfaw9A1+aaK
p+bzI1dTXfnGEeAT4u/DG9Jutxtq0IMElS1vNLwHUUzEO1zKZApJLsplQzmgAGgfZdhijp/ZAxCf
oBLFqr8dQTj/XrkxCukIcS7e798h7HFM4gZ3ZQhzulh0Jsnh4yXnRK12SOYJzbb5MFEpWxTIrzEG
H/51qNY4lyIbv+zSdUIZaZ1E0ohJVWXjTQEpHBwUrdmXZg/GRNA4OQcb6EvGYQEVubcBwTHkz1Ot
qWakZguwoVagHheCy3xfiuUvCzef8IxhAsouMlkvJ6AzL7JjqClfGWT+bkGhAMSrUV1d6u3k4ZBi
Kj+YZg7PdOeo1WW/syNs8G4rNasRDU2X4RjzTT0DWI5SXGbeAO3+F+TFRQfjMpyiyh2jNMXbymZS
x0YMjJbeJP0ID1yttTwKK0tTBPp9Qrvua6PBHxp1XM5LcpWiBY3O8MavemyC7aYexImr/IyUhhqs
1tgBFp5KeOCegj6/Jmd96CWg4OCAmNPDIKuCXLTCIsjhhl2DoxDS5TxCftzwk2C+N2pbx/ZKi007
EtXRfOxaIu+tZEWE+Ch8eqx9PGEGJ++hA3llD4r5sHM0UfxdAal6wqxaYpLOZqYp7Gh3NY4wUuAN
c7mzW8Ah5lsWLPGm3eqLlWSyGeQYS5ckPTfSCPJq8ftOchPNYEDME6yadIPufU6blsMTDiiybk0j
vdQtxb22s/mfB5I0yBc3hg0jJVQYh3N8Wb1vhQBaAySyhWkcuVy68TC9WRdTjrkvkYLNmBQBQJ9g
Zg/CsRpLqjEABi3n6mkItoZB9DrFU9YBLiawUjb2ENgpLflPHrMuktmtzpOhq3fn2SegHlE+ukfM
Oo7hyLnfTaXSmlRRqanImCY2ZYmJ1GAdy3JZkUUQfIVCHcL06TR0yOu66XaJOO4m1DKZxdB4S2sw
HUarfXLRn7+y1n1v9V4pkD319uyTRiWaPbpN6l5Qt6nzO2VeoTq8oe1scWN/4C6yFp/fZjQYayBP
EF3CrgGHZmjJmPLXUOfKXIqdGwPlFE2Q9DSw3MoMIARcrupsa5RZk4p2IT4s4Q2Gt5PTZq0cfr3G
IG8+9OCHEssOrjk/hCcl/SJqQOMif6SVJScEUafmgzvGoEpSyeGkL9zmxmTFbR1g5p40K8AYVW4j
/vWP2d4jA/Y+j0XFMNWvwsWqk0xeKU/MbMnrLYMfqf6LBAcih9FgzGo56lDJTxpdTonWYUJuMLPl
6pQnbjCDQmE80znTu1dY8cGx3VqZn9LhUi83VyIcOW8I0Yx2Kl2Bp8itjSoj9LX/vw4nD5Wbudsy
1SHhEFN5WoVrbzP+TVkjNfackQ6MIs1Bz3MRc67L3ZxsZDFD0nZ+ouogO6z201+2y33yXoWMNsmu
CgyA7qY+dcsU4xo90nk5puYP0ceq8TcXe0nPGjf/i3qrsumX0TadwvuSosLr0KFAORcGXlFb/UK0
upkIKXvz6jt/ETm7M5gdGte0L9WwMULev+33wZ+ODfi/yfqVKcumqM+IMP5/BwBc1mamaC2t73Qv
AS2MvYjbWZ6jKB+SHShYyBgbPtyn2jAQ9JRCiz27Ok6W8FfryO02jy4qh6OwQEvjI0KV6U6/Z8Ht
ImtyBy0Ofal8ekM1QFwRz2mWOcV28QXw7ieIsKWmpbfs8Dh+PwRT8d1q2sl04Jtoat6J28D0FXa3
rEfci3JfebV05IkpPjlfdIVXmO/vKRNyiuETeTgvAi6yoQB8jchn7zzALBe6PV7rU4AVfthVlhME
9kJ2tee0O/vCmzIRFt8P2JmnMtz0m2mGJ3nh5PHrQJ/6m2znOT0V0yiZ+syoR+D0+PN+4F1wXhTw
2ftJ4Va0rpuewsGJ33qVDK3KNbh830b1/3RZ43V+9dldcRwKHC1EqD0zvoa8lV/s3CFbpZIgkiPo
mNkxYBmHedBOek3YFgJJ58JBepjBusHfCNrEzv3gFrNHAPRSq5kDX5bJG0vqbR0NTpNgzTtsEWGZ
QuUUfnJHcxDPPZq9NzuRqZFMvSU/rD+8HyqRnnmCj8a1fRxkAQXoVKrFilOegAS6jPa9aimv2rgo
RuDRgc39yZH4bhfh3Gwg+yBa9FLYGKS9UO14dBKyKKvnjYWRmsNr5gaiN/DUBcc+rfyDGsdGr/+P
YyIERtzJ7hUVpD5TTyU2TwEpOJ4c+FDQJOU76Y/kaY3kA5bfRZhrbCibdm+pE2lzrldG97rujF2d
gKOMY0ayEKRxk0qFeVdnv1MvJwh0Qqt4X3qGaB9BQhvv8o1acIBSEWUtk8s8aN6u+S3S8Gr+3PFL
nSLVeUG+XPQlZVV9DJa4Z6c0HNmPdW9u1ci5DCuvhboF6YJiN87DCafkwFDvaQKvZmQDbsQjs9Il
/UJjYGSSHmhUpP0ik8Ev/vTyd32yGUsf7zXxmGffc6cYyaMDbxMCF1xhS50bRbfoV8RoXyND6As5
E5uWpnKg2yj+PRACK0hmpCoAZdDVkjTAc5+QQvVv1wPVLAgP0nRLcIKBgDkgdwVb8BH+6DDW8DIP
TfAZfg5k2doCXvzcqc56Q+AzxglZyeRn0DJSVNo81JfP7sksPQkQEdYAC7uf/7UkkmqLBYFrZWaV
Q2tcy4bxqYcD7a+RNYi8KO8yc44LNmgmVEcRmLFcnp/SVZjJl8+4o8mA4lhH3F+FBd52iolUr2N/
5T3Y7jyL5Y7tPq/VR75dvuvxXtWu1w+q4C5hc4Wq9sDPz5NvOWHxhJVnIu9Hx8o5/djbBjonYRz5
MbcSi3fcVcQwRWFkcAgSC927SthCZRtHbtB4e0dBVsDNwr4Kw0TvkW0Abwg5BJPDmD/aBrbne99g
pXcKMuNWw54QkI0X9UWH0PFSbaIaXFwtiY+mGX1otH1p0j7aD8nQ7yTXKkWcqmJJ+fCcN5BDycEA
B+FWiq5f0nqGumichW/jpxfOmkllxonRT/beKRXbNCd7bu1sW66yoS0F5giDexKJAB5Em9Jb5r7Y
L/cd5vU2XbtBbrpT2uo/XD34eboVHqpp9V2k5+VE+4xZwLqczFAU+AxkojAwaG6TwdalFYMTXA+2
ARmGq2ib0YifTBjwR6dDB2dofofximRcQ8fUK1pPcI/QinF4Rc3zhEwSe/89iEneRtXfg8QlLIIQ
bv1l3Fza/jFYQVG/g/DNiyCTbRkxrcSOmhZkT1jS9UOMONOX243rgwGtevBYgaHFdcfZBXZPIoId
3tLiJ1GHVgEHtzLVm/D+gKaRcE0t5KTSjVmmsE64dEccz73NjNXEjsBTvly+wWFjFWf7Kw/kw4wg
1wfDpf5HbsplYumHoATj1uNV2NBHugC2hJJESmhk4QLl6bkQNa+pTzv6SxLu/LxdzBsUdwyScRZa
DCiWXqavap+13Y6beINomEMsgZ9cLX2gJrp7g0cHArVt1Gpg6ycU5rtzwZ0EuQVNWrBKr9Azlhi1
Nqe2NCgt8emSr2OBdxYvC7N9gmAjNC/4malSz5y87q4SEPnCENjIbl2C3xx04zsww/kVLvEMwgT7
arlHPPLn/ZH1YTss9pzX5N0hYM6ckhQeLF81FXrceMnppP9HhC0P3QJYoe/NTYJ5bRy+cF7kon4A
grSkKm7n8RNbjgmZENCi3Y2150TvW+TcDsw39PYxCTtt6WUPJcCLdVSBRYieIMwTXyRLtCNnCF0/
Z+KJhSocRFOZ4ExZqokqEcXUZhv1zVM6XoKoALd9T7niqPwjT9TaFFfgBRc9UO7lNdt8+MvikjDr
uv5OK9AU7dTDGEZjt3QE2awf6QFhghH1jZqnaXLgAz6QeB3WraOdI3YvAVHmp+STpMoE6a7LawvD
e3lwl4A26cpoZspMLs3ErwZ94SeRSBqQ/mpT04oVrjfF+TU3xalo0ce9bwKbGfLXLxFyvPmauFVj
T15oyASr9JO6PLpHZDH2VhOdBvSuL/L+zBV4YnJFA1HBANuh85K1KUxI97VDle71j5Fd8n8xbknB
WBy8bT9I4CWggv0E8pUUqKEUtANux1kcPaOZJ352Y+jkaORDpgk5DnAlzACEUBTG0IC0qtm4/pHG
5rggb1dISmjX2DOFaDK/uVdgUaMHIVFEpgFunKaQCsG5j1ONU2WFMq2IR6tQhHpSswiWnDJOxT63
o6JU6pu/HDJF+Q5IYvU+WYC1rKu+3qJFa5K608ih9wIivX46egs7N96SHSNXKAtsZMCxonGO/DuF
+v6m0TM8Sg6YlCZyYUlcXHjRSb3lKfUEdn75L5sWb+G+cAJhJvRTW93kpZZkjHUEO6xvGqLRMRMb
Z5GDVZW62r5FJZQoDm35d9C40JZ/PY8AadhXgqtP6BUwluFscXq49cnbKJZPZI0dh41euLsxfPq8
cswt+tguJaaYyn3TTakaEf77OyBlDwDvtuIMgLsYWf1DhMgX58JXZVbWdepHAX6B6++VZ7+Spnk6
hGZK6pxGgZq8+QVgWjvKGP5IBXoQsnvqXviRY4HqWMbXeRTyxRY3SYY5nuajEQODr0cUUlUO603s
RylkMJ0hmnx9TlcAvysfeFtCxlreJxpnfpBIpcpPiAa56oK09Wr3cPcHdGw1y2N69aP7utzhuczx
bqVXg3SREtawNngP5LE+8JAmdIFh381dA3Zzy272YvxcUFWuno4Wcw7L1Yvn4ASJTIn+6pYyJGLj
doUK3AWrdo8KO3uoSB69uCoaJx+sWeM7eAyoFfq2O9dYZkzjvsrMs5ahKaJ3pDzKu1PrDzMlwZaw
EMIOEgauOHxTcatB18IsmFsqCBJByS/7iajY0bEy0RfZrOU4Wgske8kA17+SVNYQTEdKyfbS9ARr
xVD3tXWLTGKm7GcnBfmPPJMj4exv3bQ+KaTRjJvokT5ijSyn2jF1ZAsJzABo8PHhvb9q8Vh8rHWh
a/wrTFqUXcuVJLr0ZitbMstmSPTUW901RYGQM/JyrxRM+VbwbhS3tPv2oQ9/mu3rxpfIHp+G85Ee
dZ6Be78A5Vs5yCWXgOQ8zquCBtkDDSGStioIjVfsmFNf2qCbopsJ9bJNWMLiBgfWf4QamSH6HVX0
rt+eIONudvwxs80D1UKrCP/CJJXbHSLdmnHdNSs7/Kvonanmf/CvIex6SKpNckSv0uUeguaaHfiC
acI6UE4hPEyJJnjgYAxMrG8u3jpwqtlqd+d0tZlFHlXA0HJTFGtceaj/yW+i8hxUmD+w/zrFYfG6
gU5iGWBMTZkTZTTfVN3v0zahNk1r85uSlNcNNPE+NV3dTL5NrUO/f2wti8j394bTKQUGwvOl9swp
YyS4j4SwUa85UpWKL6CTyOcFMblXoxEntaZ9FFP/wNa3rxvoYOY1rlJMhOKO6tNE98SoYGcVjB6h
FIxi+KOwYUbjMvE+W7qEhNUZ3gJacP0Hddzp++UJBeUwiRzPFAATDGL/LBoByvkcyzpjaBpZvNIG
3rTsNwWHTOZzEMOVWgEuQ+LJhACi50FHRIxh5MpZYsWLmyAs9rdl4iyZsGhhGwIk3dLJq2rdfaYJ
J1YiAm4iYpI086kEZtNGgm77DqBPB2q/5pKn28phnHtSBY86auzmVIN4NzIMHLlFDrBKlQ9/KAHw
tiKDmlbDgi9Jo2Ei7FRdg9cVg7pqPtNfmyc0i6J8GI0LBYhZ5fPD0M2qj1n3Fbalycr//l9OURz3
jkKDZK49iTV/csZBWM3fDRcOjE4W0q4YYm+rKcq3aq1/3WteVvaiiRDVD5WPvtuWKmDBjxZxW1Xg
iEkyWifmQ+TdK4+k4cEKai7rgtaTSpamkPaFu+fnKhmUFz3acG5MzXCJuUQMkQ9/dMQhhdDPNc7o
ylxJIumoatOYyf1uF+cT5fg1P89M2nB9WjSDApVLZGsrDzEMhUV+dfTA87B5bL1t1GXWiR21Rg8M
g9N4xoqUVbhCARL/P7t3RYkvOW+YAWR6J6c6jKBVmHPzjbTELD9qsk2zyJQ20H59aZGQFqJLV14C
FUcLwQtgV8mYk0CfNGm8ZNDNTuACjrW+a8aWoK0M8hIUXPMIxSeH1Wz5D266KRqBhWFtKU5JRfRJ
AnuF8nE4+X/GdomS79jxmt/PByJh1LKR/PsguFdDUZpa/o/tpNEqfYnFbPMQ806WFS3eA98knxFh
IUiX+u3dV6GP7yAcCndAPyAf4XbGRAlGYdt61pYpuf7u5jajlCO675vSLeobGZfUsCWZxDHb9Iws
+lPdNAFloD+a3DopqXAKfokOmaDsvmBPCWb1b3AQeALOCTSgxi//EjUo8it41By1JgqYwkGR5m9e
m13Ptb60XlM8CJDpw23NBygkp190008edsNpNGwS4lHLKGgbODSLBPxtBc5vLPirfmvkodqotIFC
XChIu/RfI6XmxMqoai6aJQCjgmZqVQxqmD/jrnaJhc4Y/pMWw7BvowYoY9i68Ps+1nZE3WQv5gmG
tJ/J2bwohjCOKok5w+EI4QV/2aTky2mLlXD6LflKFtGvVZCFtjlwwJ9taEEv4iSLh/erL7F3ayX8
nSxL4/aLtuNJu7Ggi/xzI25fAdq8j77qgz6K6uqMRKrXI3F6AUTpXiAEoSvZ4BaUW2mcaurFm0L0
pVtnfZAHXeAN23O9I+odrl88MFTpQyd9z/NZAfWfsNG2XEGQ254pNwCXP53S3MzonZr16lJaNCQO
7P7dbXqhx3Ozs8IjAI7mkbLCYQ80GLemWxdRJgBojLdoGopS4ozSpPOHGvKetP6O8JD+aCargrf4
xfbDnnK3JlAjMFp0FZYmu+kPvOv3juT3sNBZAyH1phae8+/gUd5hEoieQmAOUuSly877PWC/f0B9
iEbARC+yIchYucXB0gvQKICBJseexi7eRN3MQkTvbqmuPgX+AmtKtgKuyv/4a3A9Gr7PJy6igBlc
Cj3SVWxBhIeQhcEZNgxzzcScBqGxGmektsA1wQM1qAlq3wSVB2mz63qpTj7C0R2rQCxwvqiST4L/
xkrxgV5HPEwqrRZP0xdtS16yvp3ZYG7ooRai7T/wy4Pg9RVxGPXTFTjJIuiis8EEK4QizWVARwkY
VkwSY8XaQQaQysnfPt2gmL9tRpXNkbqE5W6MJQPtSf8HGCqOK/C224oqaXTyiQ2DNCLRz0tPEsvw
vAH3zVNkqpT62NbPc+reQTYOYzxvNO4ClMKDXbLZKz6ThVx22pPS6rG/t3QrZq0j1Tm4mVsgxU0r
n2qZ/1pVWlmShyfJnfqYbzBcLI17BEDXM439rsHkMQhji+6M9uDYbOhfFs00PHjsVs51OBwlow0N
JrVxD7jyGc7zQ4BiSxHpbwtQtcY7dxh8M0OoxXV6gB0FHkYbtyw02GsbqExI6/D8Z0/KK7xNePYm
DTKBDi5n4uN0Pl+S92XsX6a2GewJpBhC7CxTO0+lhdL0cPerxM7rNU0Qwn0srQUt+HjwjLqbHJXJ
VB0rKyfO7XMXixoKckZ1jmNoxgf5D9kcvaygPTwEMWkAoZZhzpGjHmykez22lJyNNTI5whjcQL0R
3YtG8JUbM7DBfUj7VHlyv7kbIs9BCveO4N9e/PKhIiWFwEYZzjRLtQ7yX9aZ49TUr0c4AGa/82ph
FmykwngoK/4OCRdJtjwUt5pLJeVLYnn0A8uNuBcBnn6z1+a1vhzhlVNIlFcgrlQOZI/DG/7bRYf4
n7D2rYMQQzeIezDdTqp+KAMbxWtNjYeyvHvRE80VQX76Mq9WCdizvlB/bvbenwCdbMPjO5J/JoFo
uvYrI0hgssKem+f2BWIgbz9j2xf6Kh3QbpAGrte2MnJbpqwuJfDDwaoJWnIz+0TXCevetPLhOMU4
kLlDkmmV60JxuCrucXHp8scH6SKiZGKRMkuVd4jZvboPAnPL8f2Rz2DMTgXn5qct1Bklqrm99gW+
uoN9sPx2HbYeNvE6ZXm09M07jSP3p7uJD1MfruOkPB9uPzr0N0xrDAHb6ABrtrA70Hy90u6ZlmjV
rxvXf8SYocR+/4dNI6DGLXplSZzEYmcOgO7R9bkSvsb5UtrDT23f3RqmHlA5qn+mWA3s3sHQhhTw
aEe12qbh3/4jpUFc5YSY7BQbP9UonOyeemzC3xLyBqeePttsGZgx1K2hPXiQn1ivRp86XGHEm7Ns
rzhiSeOW+75PUeBfjNcbcfMm+hFC28WfN4q2w914nMibK9a3BaYDQ68pimQjjwAgPD/jXcUPPkjH
ma5CtTSKSdhP8Vb/9+gUmJoxpH+QnQQ1ZjH7ciltI2GJS9+Sd+AAVDL8zwKqY9lN7xPMOD8akHY7
aVQ6UWg4hxIDrL1cIs8hGT6i6RO1+nDiadq8bERiqTdGDFQGZsYWgD1EvfFmEMjSnsV/eCp1ILEn
uPyfYZ8LANgXM7HuqW5S1t5TWXjD7GtVXmjblZKEOKT6AauUGtq7JXKsn/QmV6JQLxMgQRvIRm0A
prZCVYO7OEizXI1WSx8YLNePFOkq3wXIRRW6ewKuSkUtTcxni/h2PF+0PYTU/8Mfxr3twFkYcDHU
Hhyi6exLSnP5hO2su/kqE/AcNpwi2l9Q7xlS5v5QVIDL68IoJzqkP6MWZ28NI1/As+yuhhZRZXdd
R8Esttsz/4BMedCjU+LBMMsB1o4Nl117C2D7MND30kO5zMfC1zUNjZx2IrRuSOkUWFnEUw6RGqM7
5toNNh/KyLJKTBZaQgomr0iw7kaofMTwXtds2FEi0nDW5MvcpFCRN1r2paWobDt3UvOD97YEr3/y
3w3mBWzB9lJ0JL2fXwPnRoYLURP+RtE1ODEnHAOt3D8WVAbd7aV+ciU+2DGjW+km67qaON6fvf4q
62i7AJJSiUeBfV305okEnQvu2UjBPpNYYEXeBH0eaLqx1P/vSPX0og+o8RVwtg76nXWqxfmHdmGf
2RVCAQa7+J5uMJkPwQ5agVvErVydxK/hI5zYz6XINFZU3Nq5Ag62O/bdyalh1sX5HTCl464GJ8rG
a8+caxj1mCt91NNLmM+/nrUaE8VJoqcv6BbgYiCFY7l2SlV73IlMDSeL2oKfhrTPznYgq8c4EbF6
oHBOrTlcXnIZnga2A3qQzCsI06A6mCYON/Y7Yx1gHdHvBSb2v7L9BM2lSoaYgjxqXJV6XzuufyPN
qA3bjN6aSLnYaiP9PcosKIK1oVj1IIaWK1noSDhvkUQIEa5073vTT6UHkZpMhv5Jfgyrl3vUIFq9
gYRpP5YnOhDBdAqEULv17uiJQMPlXvRGMgq/LGSo+XdUvNe/Sm72jIqJ57GxgxUW6YUmZJmSMpSr
9rtYs7iY2JuIbg2gIb63CFC/BDGxaSOUvS6mR4qSeM3W/ZgReadAnxbkLHKTNn2lHSU3EZ+EMwQ8
dnzYl9MWnRO4W2qY88qpuUHYwxqT04MMlTgdTVnFVkMsCJ85Ce4nQ0SomZ7hzAfCOdKVwr4ktQlG
hO1JT0uI0fO09Gmj8WZmkmCWF8o2AraTJEgzx7ZtJz4Q2Z/BepD9UKVTKUfqVsgOadunZ3zSukeq
z/lRWqng5Gh4G+ZsqYytSn7NwfP4dvYPNm/hNk+E6NvtTztUAQaDyT0JEI62HOKUGAIm5qLQ68CU
RshcYNXcE6majYnQyZsoc5f2sZMwGrd0PlQbwdEf+e2q6u0S5BsCUVtwIst4Ing8ZqJtl4kijt+Z
mV+dKQxCy+heZv/7UkLtWX+ZRfDft4b1SgI+UHJ4iedwP6f/aBbcX5iX5AoiuYQpMSIhnoThOG5n
4BnbYcleKZ+Z1jA0vmntIFUT9hIi1djQdpVQDA9Y2oW83U5Yz4X830zl/EnXbOYXU4ImRUtby8kd
XxMSaKS7h6Y/5E9H3CdOgb7H7c5zGjNhy7NKdY2k09mut2vY+BdQuBLJlfRzfjX0eYEveNaYHJHG
6egmXd0Mi7qWWDzbwoufziHOQDAB1+9CgCGHwVeryNQBKeaJV6mA7dCoD9yssPc65Kp+fQ565Ax4
VW/nCyT/QLcGskRnmpf3HM5V/EHlLmkZtEQZgRSZgcbhTTFeRQ5ma1cMychHnHMLybOKSs96cZYq
MRyMTlAKrKTTAkwH1+N6VVQ2OD3iFo5xzqfoQKCnXomdxFTOpy9ytg6O+iPFWw9RGjPLCY7BvQxP
zD728aTEur15AjarqYFOZ7Zjo3qppT1zKvctlvYO3qL20Gaivz9ZCAb7N9u8A8RXEdo2sjnUzoTl
FkCTAhDaOSaAb9XSlMIkCeTZ1Xl6tq73XGue4iMeqcFJkk7qkm1Ew52Pzurx8rK4q2ZMMhtJXZv1
39kuAZFCVKmlXxjnJk3b8ml1WfvGkOGd6b6uWc50QGmy77pnQEhBXWWIM+RZnCS2NxL9+7tTaAJr
3MHTeQKVd0uK42byDmYEgtF0M2V3gvpS9ykBAwG07IXfppJR/DK0QzoVJA2/vpHMmeCI5gm66hW4
5Lx2hfffYO7CAfiMxQQ/86L7z0BEit7lVSvSd8pMn5+EVVG1uPLuI+sn4Tr8TDEDl9ULOsHGbwN7
hWKwWp6EQYL6J9h8ggsqodd15UafQCSp8ex0eKzyBrvLEMUrNvPGZnSdiDnQ+2bWQf+D3nVM01zM
x0/D+16fQrUsDew9RRmc/75x3MXpgJdNTEP71xYg4QaV5S+A/kSUtFlJcZCNFDap+ax98jFc6UFp
rKgmuC1AEOa4hHvZK4zmGYStg6HryMOZv+3igFJbIzUUc062wWY8h796pGRvmmL3gb6xXZ/4Hxiz
zovlRx7QKLV/VjR80BYB8gvW8dIf2gl8CU3mSHeRmguNcyqognG9/nP1ALM263G7JW/XGIopl8uV
Tt8Crg8ugGwqEy3V8oxf/QquaY2Yuj1qobBXy27lT1Qw89pQY7QgiNl9a/QVOWBqdtyuxl3v6sx3
+avOfoLCbBVy4AydC+hzF7q3y+y5IFYFiOJ3bD/Ii9KmTJ2jbzdEn4ryso3Zt3gLmA0sFzAQ8lox
StopkcK6f6c2pCG6xZXmS6s+X0XQHS9F/n7CszvK9jJ5y2k4Dkpcvxv7SIWG0UY+N9c+cZnFOpp8
wEeOESSHh4zEtCCeltlfrnBqdznBJ2CZVbdLORmk75PuxrIucUj81g1i7gAT2dmJw6X+FdMgJUPu
cEfK3OrtVXo3iiqF3rMX9GJCzRv0ud3oMyYbMtw0ajn6ykdfnhSXOdpPl2Tb7fdhDFmT/cIiyEbQ
Nkr6DtExeCVlrKjZuP1gonow3vFPTsFSS95lNiCf+Jr+hefnNqmdc7QYx7dv/ExNsJoJxGhHMmp3
oYJvUXBuED/1ir8NgQ/9SSLjR6GKUyngkWMU/9tH7jSUhXOmZ1dQ/d+QKZYUvEjLarGM0gjyIGtH
CEzqzTTq8DuE1LUffwMMkgVUhqKaVWGowCXq4iLnRLGqjEiQAQxsq0jtASqEDQonQsef/oKSggpl
UXugpVm/OeAAR5YH/Y3vA3E7QbJUHuHnxnyEW/9t9CxTgQ10UnMtjwOvvYsXkjUV+rTqTnx5sOe3
6t3VgcSqxvD3zQF+TSqHBRSw6I5HwvAZmXWjqT1XOWUm769m0NXMdpRIzMMUEkZt8q68Wo2rI+uW
UZP4uOggeih5fq3HALkhnYpv3PSVOUb6Ul1g/iaIFFCYz+d1tY4C6V05dYXazmHUqzbFGz2lW7KO
UrGGgDBVxHuU6Du4j3MLt1QXBeStVmQnlsKWESDqOFEawigiCJVlcVEakl2fd83ScgtyHVz5G1qF
tFmd9SUY4bzP2E2stqlJRbYRC/1OVnQVfPmVRmu58JDVBNOLckl38KUH5yqezvoxxIuM1RTMSnXm
m64FdRWZ4YisrfKNo2B34tMBFIO+Hu0ItaKJLG0LVH1fbxjOonKzozOBOBNH7FyOUXbShPOXuScR
IuUNIwXwZARAPC4ZvxgFLLcdgSnsaVT8GdEx1XBzN0psH4J9gsBltAA+RLC1pNvBDaa3EPASrkTC
qhLcsUJjnRwH+XrzclKeLSemBHjhj8qfwhGpjAhtXc3aeGfd19dBKSIY+bGHJB57/fZjBMlx21Iy
cpJWvYCswmgvDrZ8F+B6ZFSMvEemNmegPqDv6YYhC84okN6spo0nVLMP3Z3uuo2QtJBTTH0GBdki
R97wTM9Uqn1XEMNEz9/G40ctLNKRBiSMWp+Z8sGPv6A20u556dfIJTdMvc7oVcQsys+2S4g8dKaB
kzwar7++sZ0ai20vTKXBb8DLh+sLn0lsOIEjN/3YuJSqZs8Iy2JJhpS9LnuGF8HHFy/PEW8GG3Ix
ylpZn8mJc/5meeyLDEwRdbtBzoeBoq2XeD4sQ1VHCCm4Yf3/vCxw+vlqJvk7IxGBWUsbyyh5c2X+
bWG8kty5qWV+xU6SQD+K2JVb6m1OWbUXDSYF1lknOtms6g062+2LlM4QJzuMvnedMIRsCsv7WDG3
ir6/tl39wDru0TZhsNKvZeUBvxb1hdde9LTxVZ3AtXAJ/m5gy0rjzSS3OJRaK+SBaiQ/SQpEw+AQ
1IxRokSZutpMwA/jY7HSzjjCOYgOK42QptZwwoB0bdFSvvEP0xYGvtUgb7Nli+CekD1fFd+F5Vmc
4hCJbGvGeyWRSzuwp9GPgwgDxKB5oOADri8HvbOPb3g/b30oLZpZLV7LWmKBjj59fZsc2N38Q6VD
EwcFHDvTTkVJ4zYImQ1N/8l9fblAUvbiWGbmhw5LW9ODCmVzxBAq0chH+dEJO9hwapzrQdB5n6JB
vbBuTTRNZ3DFqnsubArFO4LHHSFFvo+GWkK6xEoo5cPDk9VqH2KWnd5yQM+4FgTJ4C1hsvMhD3sM
CP5FZa43Uv8QXSw0Oqxo9aG0tJvzx5IWWqL6A/o9Nr3RcrSHB7dgheTPwMTHTji/LXNXbwJWdBib
zYt9Wsri61HCNNsqtH1Dm26jJYXLz4LuyFYjw4p889efefQ2auoMyKSkepqlUBrOGQhnMc422JWX
exP99fioo2eojZ6uy59pjLyTYuLX8Z+LnYTyMm16AeyIg3bZlTA2URZznsAreCcz2p5wtXimdiOl
s1jyHIbPhcZ/aEGnJA+t3dqwh+8HPja9FX4TPmbOB5uW4UQiK2Sp+iVmqO5c0qPJ4hW6pnWPuioZ
h2sczCMwn3U4unaUpyE6pqLhWv4EFfpMzCC7gxVy7fE8AM08y/aTE7hb/oPTu5jeFHoBn9rhJFml
6HBLfG0dImRofVrSdrJlRrHdl0cPIfb+e7aI44sn/dpOuk2YciyeFBCdm3wAjbrBNCyztdIwz09P
43orK9btHIjvO5uoH0FPI2nUs2ceyIL0DdlUXCq+Brsm6gZlcX0BElXmpYhJuVWzJaA/oKMUICqY
Nfnnfd/EYaQ30ofTZZAKGjPKN/ScD6CEaKfBQ1kh6N3mkuZMNKUm7ug9J+m3ibdXEq9GWqPLt2an
bTyNXk/CwZcp/A30TiptZdUFiC4BIA5kGJn5NbZIEDS8Fyelz4LisPMOcQb8x5r1bmcAt8rrgizW
vac469I94TSzz0KNIgW8kqsHgv2vE5VQem0sicWITC0gv/vIFdYmhyqsL3XlL5pIyPCNQRx2CrcH
LciWvUwO8sfcfsWhbn52MlycHfAUXeMBGsXAb32dv2xTaYP0jiWyY+6M9xeJwzo1lFqjVog4CD0C
gQSHAjhi29HNITAo6jq4vIT5nXgB5U3/KgcQbWhCrzzQU0AOoLnZtNR8Bp+oWfoKaS8omxyjqg0P
vd/exzF4kNd0jVO5ueSu2tEYHKz5y8Htl6OvJbJoR7vE7C1D/+F7aQ/xEQiN4sK8mkT4Ew8N09kM
k3hpzyT7VwLdTrXMGTorEjJnWnIXau035XxihjuQATdBJzW9wQqt3mAmSTYyNF/LYkcoy4ry0CCt
mVYCNEpR72Z+vTS8J6bVKqLrsEFUxWnBuH+lvP1u6PhC2bpxukccOxyQUc6dwIwit5MSc1YFEdR/
EqFtKtly7JoHzvSuFndrFrm7WpTBrzPf6s4GJSyxX1a4iNuGJdvynWzHACcKLfBv4k78bTdSs4cp
MHl8j6ai3mg8p+A3YCLGEo4Yu1yQy9m2edB6EAEd6xvtH22i96SOQRVqGjiKy4Axou8qDS+ClzOf
msuLXtPudndgNBDRYD7RgSPiRTEr81ci395QRIMKdQ8dRWuF1x31siVSpOYGHi4M41993Yj8M0+D
aQbljxIkH0X92Bp3UxzEsTgCROp8kjso6QdvB9uONutov1Unz5VS7Yiy7UD5EN4OwHsTaAWnjJwT
qwdkLJ7VP+TEqekHXXh5Tid8JUV74SUZXTQ6o+QH4hGoCn21WOT83UIW2dM2DriUKLSsGkzZxxjM
XI+DDYA5aWki9X3yPm+9vQMoHvJhQJi0Q+j02ELywr2es11SWCaFSTFXH3sqcEuLZPLXHY17wEoH
s1LB+USx5WcUc7rC2N/7pb5ktC+Bv/fyveHuVamlTw+pGW3FLRWd7Wxn3A0dByy6uQdwtHHIP1BT
Vl1o3qLd1+S3KvSC7C/YR1hX5GZ7INmTsL9jY2PIwaIH7iAkW0VWDavWOj6IaGf5HjtskvXN/fVd
V/8HJwNoC2sgjOZHaLEUNShDlgTjK5c060ucZDHMnyCjW2lSuJ3IQRFOH2j03SzF+uxXuZw74NM1
nfl6i9gPne5f+PS027ztiCcx07PLPewKSWHdMB4smCSCgChUTDFbWrwaMQuwgkSMEGrfhwYdAoRi
oUevzzWshG2G/Bbv8X75V+y8mj6i+lGNxx5I5nkgSm8TDQCxpyH5uGL+AvBmTjVp/arp3LFm7zy8
kUCXaL5XXtymDvOdI29d7tHr00KVr3B6Xh+qhj/6DC48NmFX/Lm+UT0za5wIi26s0oOIi3bGWUT2
nIup/QT1hHgJyQ5t5/eVKAisvBhL8/HPaowktLcJrqCeErx1ZuQjULkHV5BlmSnelro2PRnU1gWj
Y1X3Bbqv80CiWRpsZAtvuibL3IL2EeZ6PXljbFugnzxYrLWQoH421K92+9vTTS7uGu+wgEbx4S+Y
lY/7AgOQ3D3PKC/A/MeewY5ZKd0d1fRg6R6C4+K09TZ0dhg7K/+mKATkZ8Pf1ZYeytwrleC6IxD2
y7DqFwYTYJ4IWerSrLM2wnIHNLYIkvqTCrVsu+SjvakPW/CljG6fmNKEKhOE6eVFxub5HD8ovxk6
1qjOJ84rgklwRKlffDMO2P1Ic7cmL4gQi9xvrvF1XFTKgWrK385kcyLmv72pqPy+Hfmsr6qWMYnm
xRDwAedOeJwda3mzF3cpNwijq/qHUfR7LaH2y5EIODbPE5UNu8zw75xohQKpdfR0SISuIxDl5Tjl
JOZEpnuXVlEgrg4md8zt4Q/PfarnX0za5dYE7FQrsUNr0kLlbWn5UTgz/AjcyjvO0DDh4MjxpOyN
qI81VbeGqv4pyjG7TZW+2rbpvmJc9RIL99Lr+vJh0JYwOVQxk14yb1XuN2pz1wBxRCc/eu8VqMHl
iT1rAq1ZOhnwII1VsP+ojqxfOzbISROKld5YxYht8bZa4rE4om655hESXgcT1+XQBs8o9lJivx/I
xTcFqmYGnROS3fzCtjUr6ng/XN8iwvguUMvU1peVjhVXZXTriQJBaGpG8a8okYFrpp/wkC3Qfz39
Pu8vcSoVt/ct+gqWwweotMPvvGAjJaMeUkzcHgi7Urv3ORWKA8kYvMhdNg5o65BHrDaELVQXRpHM
amxW4+8oxRqi6VytCTnAOG+DWQ+TYj0bzsJ+VffZyBdO6DsNAxZsG3jGkRdSOuMAOZjp5JtPVk3e
ipVMRkBVmHUPBsYpFXp6L0bK3unuJcfqYnzHbxcYiaDOlW6trZSrZulzjCOvOIW6GZ/MKBAaBZWQ
tmGzt45VxIvXl1Ick4CvzF/qF7dkJMFwbr6thgTBM3wJs3ownsbP55aMu5PC8Wb1dZXkTD0WEPf1
ZtlyJ1E1SiPocNxmCg0lsrGLmaIW+yjP3x+lWsfiFyT4a/+KIPVJ9H/S7d+r5lSBqCSiErBqIJmZ
ttb31fsYYMWKDb9KsN6/lgxWcm2l1/m6oAvMktbt1LDxbvG7ZmU8YxidgdONayTFWC45F4c4DFec
nUURpMEfG2r7LMjNmaRCF/KeIiG/ImIKRSes39PiyTbiAbF8vBeAibkXQpMt8X3Vjop9uUJiyYCR
75Ck0r2I/+cEDc1kwppfl8lvcXI4Gq/ZwdvWFDOsYzy47UdcAVUYp3K/bp+iOYBsU1YZKhbR2owq
PnDipq3UKeDnyuLH6D8DV11lJiqbEVyCqkrnR+Gl7YgxJFLyOkHS7sFzuYVGo5vjkNnYlKeCSl1q
0H9UYyTsO4xShj60c5sIXHGIJfgIOEI7f9BINDpMquP5OrE+QKnSbcZwHZHsPDbwjPh2lZEyZqzf
EABG3/PotVKlVK1KoKh2N0PZKepwkr/y0jdbCdiBYICvp+Ri2tdefN2XFCx0DdErqfOUBfmXN35T
oy+H6BDZB+MwS32bOQampwgwwxwPeiv8S5/tdbarh0aU41NqO+6BUaFWgJkAoMwQ4ww4nBBUiSfi
8Y+lg+dgaAlp+kcZ+7X9yEwAl2vq4oH2LqdLbZy48TEwFmrXTEK3JtQm1sDsTzkdCzWGT/es10k8
G5FkyQH9prtPJwpyebBoPhU6vUES5ks31nfqnSSCIxzG9eRUqNGOYPPGypk7jlQiX+SNKWvSK3SM
oL1rMM+RZJDSRU8Prxn0f6IigL0VXirKoO6E4bWCIE3za2m0OH/HIiyEcl26u0o37w8/aQEK9A0G
kkBjf0oT+JLhLW7l64+np9peD2+iaBixEhLpJSjO2YJRssa+ALtq58Jza6g9fMB6SG268w59NzOU
ynONgBwJazAFUn4Nlk4oYjQe9BSG6mffVoQXssO8fObe0l1x6Ou/4GA3zgZFNWZ5YAyTBoSv25ql
srKyCMxDZOL5EmHcTLpLE52w1gdruGYcgRhGx0t7AS26BjI+f7evy4KWxxO+dfvOnh+6j+gX1S7u
U6clseSeFiHjIqFXDgMA72o17xi+/UQQBZu47II7Tf9BUjfmlWAgJeV5fQkPtqPSn2vtIHBpyT/M
nEIq+ZqlRtL7F6XYDZz5aX7a7RvWzpUhFRHnFJYCAUSV9lFf7Pm3aNP55GsAADx80fkfkwH2VXWQ
kHTciPrqM/6oEHy+sVHFWbLShfaRdinZJbLa0orjYwoy37Va8crXOE4jKfDbJaLuuse96XMWsCHX
W2HLPzRpvSQqaQGtK+M8w6nUksQXvYCq4KCjhJT32p+7sB/6116mPwIQQsq6U9TexHpZXqlKzA2J
OuyQ5O3tnxd+8VCZ/W0Fh3F/uqeJR27+MYVrXXUSxZAKJzTRUC0qVpAwrWir5eLFjPSp4QbA2E6E
PTwcjAJyw6jLhW9vEI2WOyrz8b4wpH5Mcx+32K0pzKNBfzkhCnuD5/JAJgXW+RbNHuvPFmaTFqVb
iPWozvfXDMEY6acIr+5lYHgzH7occ+a0YO0ZTpAkvk9FCJSx5fTEr763c0fIn5ePIxND9SccCY5O
MlytPq4ilL/kPDxb4mlNJwl195A696cRK1KiMb6ROGL/fU+ExzBiwjX+mmu9Y1a0ukYr5JvZFAVz
oyjDXbG+oHXvtZ2Wyl0r1PmzjddaYXKONUWxanp563be6S1XIGwvZieFuSslBXh8ZtVTyACNbapg
eQ33IWGGAGKY7oimsuhgOxBvio2MKb86wNCDZQTykSrKHcuFu7aiH4VIdz6juPphtoSaC5JqNJ52
Z+gxK+04X3xShVg0BU8LYQy5fBPZjoy3UiJTO+xqqaD/cLQIU7lPYuNzDIes60Nd9k8/utameRIj
cEMLpfXFjTiczJOjV50ohDVnEI7ZBe99wer8/qYafQg0xPm5noefKx2H1E2oSO8U2aSq4taixxKA
4JEJJZA0jW6u6xIaLPBnqNcShaS6I56iPqZUr2TSGJmTHt2+ithhANsO5ob8phgK4GIWAEbfI+wI
iy/N4c2VX4+UiH6sD1dM2y3Qcijx6Lb+CzerxksEJFCxYsS+NW6TZpu3mrZ93+6rd5qrNZhBG+Sm
KffQ5mKrVdQLliwF8X0Lgpa5RjOXWcI6EA9vWfmUn2dse1mVim5f0Lcp7gwqeX0DKh88zgbBdtkQ
v/SsvdrmZDwLOb2gHn+HBIPg5fLqDvVxnIIjEPJdfueiiwxCbgMRYSxnpATAstt+YcBicPkc6JWi
f+3MD2iADl4IoVTCZYFvFvfFAjssNgNJQrP+WF1Ha4r4jV9hRWYImB0URANmXgan/yE8+m++S+Nf
YINjZHhZ/iuo8b+yaSAv3Nz4kUsnLkA909tQxwniOM9ABR9PeHGKUIRVAcRyj7RZqYaVcskdlxnc
npAxS+7CnFjV1wZgpf434Dhu6jMekQ0LOhmfEgaXR2uTdk/gmdB8s3NineEDMtza9WXzqRaRWeEF
/YEI3UaBfT16q6M2bwlyy4/lA8l1I5X2rAMrkJtwCnQKekrgL8K45NfJqv50XN+37eUjnRyF3TF+
50KP9owh58K90iRs3H99y0+puUQmEAOIN3HyvrBztMKJHNQ+FqNV21W+7SwoJLY99LOcPgCJlRo2
Eh5Tu8IM+ULMN7YLqv7KhOagSp4jPaCszHvSnrE6xS1W2vhYy9Oj70g6UmWEb6tG/UD2VPWBMI8l
YeEQ0PqgcyJ0RbNcB91/57/ZQPYR+5yPXZtivVvnhxyOJCzx2d2wLcvHVluymYzbH6eaB1q4pFhP
fJC8V2oJInBflVCjzC08kpQ3OwnZ8jgMVERV2EnaMr5vg36e3nbbDO0q7aI0+Asn5TfBV6UP6zzh
ufXuRc4EjLjDTMxV2J8OfWmsWcL+5sifZcGGXG3Vk8M/beGbaRG+EjzuEGsNF0R5e4CsytGJTH3p
AZcXLgUp0iU2ws2ueacpsbPhunRdg9Qo58wxJFaDHA/oB3dFQDigAbMxQzUE0ZWBQD0vXoSt1+1N
5q0EakMgot9/G8WS1gfT/gLXmjIE6QSgYwS4WoPwBYscFajpG00thZrwG2jW63R0Dv+6rksd7vzf
8agje8aV7ifucdqC41NS/T6kXl+yBnXbxbs33NoNYNuPpHLH9E/vP7DVUae1BHNyE9wJhaSU1GLN
9j7sHsj8onJPRSHNtUUb/HfKCsfc7vdqmmXGa8GGG3WIzvoFCKvcDwq7lM8LLHO3ho6Ghk5UdBDC
PQgsaZv6CIBRthnhepNbgM3PbpqesME3VTGXt/n1LfbzC0NZq52zDrlCYDrs0hcuk4zxEM7n/yKd
mo9YoBAeCEGsCcMkUpg95FjvxjWdqU3DiPlvPn8TXr/w+9pa5dFNzEb8zPvdtW3HM1tEDkzPZ8z4
UC6KnlSkHwpiQs+falRQEHW+fz7jOxXrl7c11+hEugVftNjMylowGNqSUYvSHFN0GhEedF6pZUoh
689qOl35H/HSoFK49likYuztRjfiGzjY3crAHJWtlnMZSbdK/ZQwoLpGXSSmSzsDyrdPa0yDqY5b
DeVzSQoCWqcGjPXAd8eplROob1dr2tmfGPMP7z9WSOZHJJzbAlPdOY/7RWSxL1E/eiPYPTXAoeJy
oul4lBImf4KmqlMmsgC3KuT/dTErauuiNuXedgckpHMzATt+Z2eRY+T5Wxc2wT5PHgUTG6GQZTGb
uZGE6e5YOz0b1+bxPtHLsRWxBQRWsKY2s7jZHI1+AMvcVYVcSBfmbKISbzVZlKvE0sgqLZEVM5Td
xEcNV0qIFnXTRO2Ek1Fxe3MvqnJJqVYg4pTLUFiwGzTMYD7cfcsXbXHITJm3WtyizTyGPeBSqj6m
W6gvdvks1UJKpbQrV9FUWtVWVZgxiiGbQ0ue4uf3aQbs5HDpCcECfISp5JBF4/mjldvoJVlwsoPC
JuJXOzSXaTLrLi8pKr70f0S2TMsGgNUMjrv3il2DyjSqUk7DMjRxtm5vUkpaH2yHJzbUzmteG5ww
CdKaXLNX+TqHuNUWNAhLNSDaM9/yKqhlTLTgU/exlHSPfgNtQ96E7FDumF1nOcsZaRy2hOn8Al9k
Kq/EwaDOBS3BGVBsLDKXO2gRIs82iAe5v/2N5Jw2wPTPpbSf9MCjVB22VrYrgYpC6rnsU6bL7au2
wQ8vXlO1AWqKdsiuIqeOke1ASs2w0ECu7MJZ2LJj9Fd0J6GSimLrtQme+61iRfmKZGW03+cAnx6O
hzfUPHifI8eLvNrwBrTf4fbC54/cLXdhpcOB5zxQ1DWB/67Zaqduw0GItdvH898tz14UxE3GK3xW
50RKBARYQtRqgHpNFbYZSh97jw4+FVymCp+b9mK7yq2DTWjDC8v1eL1qX5d/BHPgwEyPsOO2m8Rd
JgPwj/gBJ9scuUfA/FQd3FjWS21XXMJFrdQMxoFe3QGyzuNk04F8dRwvzTPH76+4wN/q6fB069dY
764EO7Or8mOlGH0UMoX6vwgkrOEN5ekxLHfxsYX0nrwZyVch7gNVmoPlKLUrgIfbh8013wTLBL1V
wwZAR9XD023U9fQhFgBHY7fr6sTtqYCrpxG1UW+rFw9vj/+/OgP6GLBsfITzy1GTf6rKLlhdKocm
lWZb827qvBHCWxjpk04ymV0m3vpsbkQBU4ycoXexLqt/KqmeijPNj+hYfef/N8g50MTxeKIeQjXh
g790afj7Vx7Cohfddh0FgH09yqW4odl5mELE87qN/wOJZDp+HuLzJcBG4mPxQUeoLFPq5DD7VaYf
+QIaPrn1t/n0i+6SwntZ0oyRuVnf/56kPk8eQCFqURMF9vvmwTfuQKty/qenIjSllBwpqGWO1x1L
xr0QN0Xb/z6Y8Frty0uTUJ1SK5lv6RPFdRrAboNuCtHhE9XTpZwzMbQG79HhF2mDno4TBNpvw9bg
p0xGRoVaAOY6wwkNppUWb/zzrEUbE0QlUfqrOZtbOjboAIHTBHEbUpukoUMDEPQoYCNhRR3QW+eG
4uivUf+9Tp8MqNOcBjr1FVFBCl/rQCjnezSmW1qwzm1fE0M4xxeH+aTI+SQdShD9VM/+ExbxzXgR
M7RMcS9bhU1CTkpRN8EJBOxSEil11LPpQTz1aQ5bKrkn43Al4Z4nNeM5UZ8QiDJG9Lb0l/pRFZXh
u7gCOox7M/sv7ku+GDgZ+xatqe0f//mMHXDtAf6jatxxplkNoNpmgeByXW0LCO9X6Xmeg4BxRFYV
3bGNmni5m3rCHvIrolLtL8RX3en8QbPLcJFt/TvuL1SROemuaxBV3K7pM/4tKxU3AJQWr+PgXeoi
7S3voDi9aMJ6xyDfxWyL+QMBSpCIPClOosyWvu3lqUqI+TFRI0Ysb5S97xrPCNYRNqkrMimzbpSV
FoRN9u9/3ZtGpkeVIDW0vDKiBFcgltJrq44nkHSUHHP2aNvtciA/agJVJeuXYHD2u5H+UFnPqiAS
kxrZhMCIZMiMgbdBXUDrSCA08pXdUZkwd/tdkgW2t5hJeCN3E4+0bdrWKDpIRIbeKVX04dPI59Gf
A8H+Xu9OefcbaB2AMwItdzNpE1UUuqpso96gw9NHDNzduccMDW5VWTRQzTGCQSy+uzuXa8aC5+XB
ZxVUU+9UOEZ2WNuzpcuCG5GAzdj9WNeovQSRftdU+LN1+zZ76V0g8wZkw9O+lKJLPjLQs+wAYLul
divWkhqDidZyGl4Ttll8WipwuuskfifWsNDXV/i2Qh1KMDq1XwPetuJRkHTJmbBjbAMmnTssNwep
ohI2KJnQmp2P0/VxY4zKxQinHIMwEoi1J9NM0F2ccbM87zIaqQEKobf6W/y/Fd046IPXCneiBTvB
sABIljxFSokNjtl+3dxPVbYDvzgeSpD8XGNq3sRkowgtE/O6NX0RfkydU+apzd3rCcquhZ58wsld
s212gYiDfR3nnBO4qRN3s/IaIL/TgM1+BVyptsxdXnhlM7VRiIeIyKUjIblc2aaufvclMIqR+w6h
WJGQmyQagLXP7K0KKl0wEIj4kZJyI/o78KjZVojVr5of2zAmiVSEATQ6ROJdZKUep0JMIilONUzR
k9Mmx1TiZc8LOW/Yndmd1GtLmMO2hxkCHK2uFAgXXieMrQEhaaA5/cZqbJYTtmrpJ05A/qhUEO3/
+it6fY3d6xon0nfeq9qvTruwElTSC5OGTUB2ZcRV7O5saukijNljm1o4ikGtedzBLXeX7FEyUn+K
gbtO7DqQzcLx0zery5u8vsz3rvYt0cVxqh7PMzzregYKaHzux2I/lkLGjPEhQ6iVeALdA9njveCh
XFyswtCOuevqkPXnj+kWUo2UrRHChDKW0rzLV2KxV/Ns7q1I/heJC+qewg8WBqSkGHeX5+QFDwFp
ynM43nv2XVQLW57bBdkAFEWOtPnu5esoDpnfZHSjpQH7eaz3Mtw6Qm9p8dDsMtgpT94dqhwmmtbb
A1CjSKiOcc4+ush9Mqp5ss5MPmOwjBGcYMN3hGbtEGuvjNueUZMuR5aVYn67iFPF8pHGPfKYVg4/
fFEyUwFLc2N4jwmM47lOzHl2ngMgShz6TmjAUl08IrJRcy+tjsPvSkTN3/jxtZkt+BH1EUmzsyJG
4eCdzYJZQFviiU052vHue896ulZ6CqciN4bKUblxuvhTXDAY0c3OeZM7aXIy7AptC08kbKiEZRzj
2XH6v0yajbIQZqEiCTYqDzS438IavG46o+1w743C+tMV4DAtQoxVALr0BaVYuqmCO0DpsmpE6S+g
MBfrhnMtSh6beS6JXUW8g8xxCp9gkFp2Hv4SEhAfZ9AcOH8PRONJLOi0MEmU51l9IVAlw1v2kKx8
tSZosEX5EEcJgAAXrYCZy9yg6RW2K9ydrFuwYAkg9MBRRLyyUl7mzZa8gEF/fLndBXz2siaFmIP9
Z0llD25MKyfjpU13xUX7MH7ememnY+1v5WZbsgSZiYTen8uvYTXAKcXvn41d5+x3YTdHV5VBLkhs
LA2o2L7Tjijj322PnZAGPGoaxH/Yl0FhKmSs+3EozS9brr7cIB6VJJgYO8Kr65QHatxfHXMCETJj
O0mVxSi+88HvAHQXS0+y7gGaFSq0A9JHTFq4WzWWRJ2QaZs7kvAS2Eqrf19pxHpLL/YyR2ewnaKq
huWUgppJRTYZ8/vk5VobLZ/fz9JCVT/4jjz4iTRljGSVPCwZe0+3KGfw7c4R4ErU8ZbN2V4bvXyd
nfvkDlsi8oEUwTgwhC98JwqAc3VcLxppZpiCR1Q3CqdADkM0UUqQApNdHsT25S/hCR4eD4uitKth
ci07nYp0crcij3y/xmah7CKbCe1kkB+V0mQyBo27Ssh9EsBunLeJEuXpM5KhaK6HSEAHlQu7ItQW
HoTLUY1fugTQwGy9HYL9qmtQO9TB8VK/CsrsT7HpdL01UOKFybohmsqgAube7+VgaeqifPYdr60M
WPYGF2jDpRszgoz1QUsYdvqVtDF3TN4zyNAUDnFbshSLr/h5bTYThxEaMoveSBobbh0RwpzvJaA4
Ry1tmEkVTICZLYTHkC9LQUUk9P7Rl0S2zmORTw7cxYZFDW4rukkayx//IesTScB+mqyz/Y/K6Dp7
x+40x2+XEcMvvN4sRwwYI90IghHdMM/5VQetpJEb88sSV56eh+85NQpzL9/Bj67Z6KxDYn19NkvC
isCJIt6QKoqE7teWe5eQ58cZ541rYuWoZyxabqq+DuB4MyBe6OhGW53snRmBbiNX9VtV4kkW2RKA
6r/YHgfy9cMVCaGL+b9xzCkT7TqIWVeel0cnPw2xhI04YqIsVMkW0tM5xQpXAiRFQ5fqLx5MoTcD
M4VYmy3XEb339RcSNxKwWpFYFZVANlhr5BSSM1TwypwMZCYqPyuytwWXw7hjmXtGjktDfc15NKSJ
kUjJniz7c1djNZhH9A+1SkqmlcSSaozB/JYSB3d76CvyFlom+vefG2WVZodUWCOrfryNGkdXDSG1
2y0brdcjHjmbl+qFdNnqixV1SXzgvYZRbE1Gby5PypX1K5CCAbHsze8qMlYMktPRXrYAq/AbEUfP
MO50IiErl3421pyeoK+pMl8rYLjZwHZM3ACtHOH/GS0M351bACamJhpH4KTk2NQRtsyEdWTHgBFR
SZZLR7DB0a5bvuFgwzpW6I9BJSAX9xvjM7f8ZYV9fyq1Q90CTIBRejMrixBQOGuMKdT99YPMDDaQ
NVzORpCd31zaxNbtLEH5n+ZUDlyfbGtKRnG3om4+kcOOEuv8aFIG/YnxVLU+V5wZC2Ig21c1SqCv
FeQlTM0DsbhCT5nrW+5BJA9VaMY7LI2WMawkq6ZZuBKpvTl/5SOwg58yiziAZWxiMrMqQ4WM7acb
YEl3dBfcrpkWNhi8PgqtHfGwqZp7g+PeWaCEebncVPjy2g8CGKdsoHhJbEPJMaXL1fX4kmTAOvqA
LMMlwtX3onW2OXWHhHUnTUBMwvl2h3S/tivxkdGt0r/2NWV5ajEtc7FOCqK3zh8cXpmxhb2XXwE8
LoANK+ULYdjUBdJKEtorCycGYzshsOdhgEecbTfQaeMKkr7sFdJ4Rhg4dlY5n7NjGK7cGFnd+F5n
46XdGpry+CmghF7jO60/vITNQusQ7eq+7E5M9gDNuEUnfTc+iwun2TckNoVojHmm81KzlyDunp3Z
wo4CzwzV0SquE2fF3HEaZbRzhUuspsjzxfLAgSAWorl9JZflTR/SZs0ecj+rsAd8y3HG2VqE9ePK
4MKFnHStIwwdHGGqiwd1/zxcckcQYbr09NR7TCTAhH3D6gw2KXv8ljUGWAA4kY7KiKX1dPwv6mMJ
XF65809LWoZFy2gNsh23RzBGjinyhUuyYFyvWfdZWobEzGz3GnLDjVPwaqcGx1lkP7VX3KQBnYgz
luifoldpWrU8gcIWABFODJ129y4DDmGg8pCztMw6qHE9PdVCAgqLbtAo2MB1ewRedy7uuFr9gDLk
XudmaJkYFCdAZ6KjXV0ZMT51rKCnn1VbgmbqmWYC8PSmhti7dJRLRFdCgdNN7LIdO/Ombnm3pdU8
tiNdqq7Sxf3lEkS4gtXH0hrQIh7inDBEAAvjKIh/0Ff5WQgVui3af07jI/XC2riBBSNIEEPHvqQl
U+ZX7RMdaTuG0GJ8jA6OPRLFNcYOmjHDb37QMCCztwUrAPDo4T5594u0ZntgkWs3dAJbe8ZgQJDp
V1iMXbT5vTDcs3QYyAKTSswVQTwfNsyB2ZaN27klhjRpZRfETszqsjplx1DtIiIPCcQw0kPQJEw/
jqZKo87usX4726PsmfvVFaZJ1LqJYktJREgHEeIj9L73xVMDBP3QQD0G0RgmvqJ7h8JIOvzBPq2U
KPEP2+bEmpunTE8hJ95j7md3xuUdPTwk2k5+GWkvGkIg44cAydN1MFGoIaTDjZf5AvzO7GUH2Ikd
d+njiw8WePG161gaN080WCSvgft+8HTJ6oajebV1ls9SOSfkyGEpBw32SQ0MMGzzGjaRcWSVxtF1
c7BlYnYGgh2n7bfTt25OV3BHbGRNccoc7hUrxmE2PPPyaGT6kl1H9y01ollwsRmYeG9rs3nKtBdC
mOkfRPczN61GbMwBZmSNNvsEdk1fkZvHnkhYNv3Kv5qbP4wh2CrJUi1coI+lDWItIo2ognPkdSiv
KmC9dqafPgkmuWlRWPjsuqMht+aH/BnvW39uufI3LGQyBmzT7ompjlgKgBfhE1UdlyVGe8HFn8+z
QzqupNRFJKg+eYEDxeGO7LTlnszfoIR8Dzg1geqFNaoPAby4zPJN48e6/KMFqAbkYOvuY0j1cf27
bLqMMceJbyK/dmKo9cIlshiUo0vz+o6ZskVprHRyKVS1fHN+JYW1ovbOHIQkztmQUe0L0KqZxiyL
AN3xS5HkgyHKbjrp3onU47nEBbM9jyNCQs2/HOX6QDMQKh5zpGaxDV88uzQEsi/YtS3aFFtTDnLd
neppWooIAzrqcNyDUVUqnGgqbmFgUU/01X5sq09NKgw/qMHje8ER2dvcrILsF4uPzMxz0Sz/6Tq+
0soZoGzBPWywLEQzRJb56vMzxIw4vN+dM7nrluY4g19vV9ck8xJbyILZ2Fhrsuice7OIgBpRUeGI
8Ht4fuvKlBvoElcMwW9Qp/VLHdCbJqAtye+kUIUE+q6akPi3c9dS8f1aY1yv0uREQvO73xVibL06
XHig4QhBa0A2eBp5TW7qJAhkRITkY3qwFeSqqDRHhFaJBr6heIwbhXZUs5gWinTf9wpmNxqrnHTQ
XaMyrVbhVBy7ZZjluPMAeEC4e90/5l0s5Biobc6B3advCybZyyZzq56SPjMmTCCsf1SQWAAHlGg6
iwFbOxtE3UO4lM08XaTeEUWokWNpjM3FGMixXZERs0J0mWR/EFV0nCSh+e7RLyrNzszcwFHqj8sC
O4qOwOidJ5CHHwo7t+Uyn2yMHPJNoe56jk56WGPmhP2mhMcYkL0PpxTEVqv6qiACFYcyjG0MxIsX
iclGIXmzc095qRJescdf+fZFP9Z20l1wQWOYQwxyQwKPG2bYANloN4iHev3EE/2IgZ4dA6PaCAHW
byusitMzMxh5jJSj2po1qAbVitS3EOUrEKvrL6CnKX78BdUANXOHhlqZSMngObDZJoCaBjfhjU4p
kCejUjodzGspX5hCuzb8nPryMkyIS7TOQaJnu+NLhfPmyVY1j54HyF+hIq/Sk/omAYwoPFMNmv3w
LYrrVnOddx5MDwumN/C1TYghTJB2dy5x/tEqO6JbWHPcJCHkmVrbW4rfFPn2e/hHvtrP0KLhYG2d
LwQdqubtFmFSWtrcsMqpdO2e803T3CrxVdA5fJGDzPzrDoYd8U3MabIJBfUz3d25RnTdFRYqwPeJ
OdIGqBsJgFG9/GWlxnVquCWOqyS+0IEW2XujmOZNACTXK7resqXgzOl6S4+RQ5qFSO1jsHBHY40j
BxJmL145ehDqGw2Ocp7UzlNhAC9WONcJqURrFL3UinO1ET5Hfuc416V2lppndpyUpYZPDZI27i+H
4Sar6UvyHEqr5IL/lRza/jFXgafSB3Q8zhXujq43GwX6MmrJp41n6AzyA51Z/Wnjft95GDuTInMa
kDLA/3H0xdgPDuVnzFtCuemkEGIvVEAGCETphPobNpr0b612V+jAV34rIqZUYpVZCfFGYpwaGLZi
qp/7nFG9RD5LttpY17M10NUKL1r/XePfVT0+6FKK6S6d5FP4Q7rLLOsShBBAyk1R3vtMdtEuXxhP
eFge1ZGU1a4vBWC50c1hlm/P/2udjzedTOlUFbLmEg0ZTip8fIBKWX2I8lRIYjynx9AokgvTEpJZ
zL998xbTiNkruQnkqGYztZXyEZYBldVuFiMEwMPIr/VbIcj0kjYP3npFXrsAkVXsf8bZfBqamgBV
GhHqT9pg6/k/Qy7tA3Dk4cHu415WWVP9w1yg87/t6BO+NC+li3qb1gGrI/67+oukd69mxY0wxZXv
4mhhL/d+fEg7DIS0mhNmrOSiXbEmwQLVcEfFWQCNgBs7WyrbGmAqXoMzEXDSzxaO4aIAoUh19HJU
aUo5t3vAc9y5JVsPI9sVAeY7dQ6EpW9SziSoQNGkV6vhYSbCp6KsvfcvApbjDBMlxlOxx4g3Att6
vrZVo87F4z4pP7aEN/P+W9QjeZEbgb7wo++87TCWPm1pvqDOYNoRS0lvvku0FwPEBLDRreouxFcX
fgGSnW3oEcKhXs4RiEsCHbatwPbjlgIZp9Sc5SPSZfvByqUxHAhZfs+SQudjhbAN4iOnwGObTxGa
dfL7ETvM4TB/x5SfT7jFQbd9eNUuiDwBI/ZzYsG+J8ShJEv9mqbqSgPCsLuDDL2nxtSIUh5OEqzC
99m3DGJ22J3HUGGqBgsCxjDtWZ2BKUdxC+VFeYxYS8dbcXldSHdObzKWV5FVV5hYL7ea857RW3Fo
A6rV5+HHqVmx1z74Vm/gkt8Xd/WEfO0KHOvCxEqFbmIg0Y6u9ZwTF/eoYTi6yYRQcBF1lIu/snk/
OMRZ4MCfpTNaO6+IujJzWgNOtlKfqZD91nIk64T/TkEmjBVyMK0kHo2I/VFA8v96+4krVvFD7Mze
9FYl4kprxzmfYbIdpXtwoVMRcFqRiygJV3vuDiXuSmJuj7mYQMaM/sZ4IfW8/nJ6QOmTrNty4b0Z
3BGdke0VCmNM+hcGuj1C70tPJ6ttH2lkfMSfX4KfCd9C+m/MU+rwcQ/b2xd6LfNt6b7kCqDTwtux
BaQbFEFc15HcfsCUw2TvhDhps2s6HqBVymMigKfnGMAV6INRyFd5Hmec4YFoF9c9d0yqaAB5coau
Mg/FvZf+G+cBK5oXDCmJPGfvpIEwqmILh3+h0K3wF8Rji15IrtGC9wEuWxVxM3rUkVTCSrLYaV4w
WNK+NpSgP00ytqT1SK8FiA59Ir+jUMLFeWefUPTKbsXugMlOYUwabQ4rXkjxK8CVSxVMiwr77v+z
g9bnzEB19a96iHC0HuExTm5RbUnMun39OO8jhwtMevijSYYHkHvhdS6uvCF29qzE5+Wkxv0Kv8ej
/wR/8kMCzi5OTnYb5naaZ6D6P+wfIj/LbPPgno/wAoC9DEwVJF6Of7ErkOKrLe92DfPhX6r8g3hy
N05Yhdjz6JPFQZ8h6ymrwmidr0IP5Z7lQd6WbxWyp5SgC9uwCyMGSGau9Nc50z7QRGGOU4lERDOX
zDvglQkfHCDEXi6Z/Dtgy+yIl1xNVWwi/mvdE21ByF9F+Fm19Q6lF/Coo2Wl6ntMuk2MYPpVvW79
dxd6Z6N7Y+6TrzotrXvUDGwObYi7nwLVXXcWI9cGvQMWJdO7vbEbcLsX3qF3VujG7AIoGVBWgnnS
XV9deSBlIxHAO38g1DiVbdkKCpbFhGaYpeud+uF7+DUdtoDMMIpWAKbj5/ulbzKKSF2iWgo1UGYq
sN1EtYrJYYx/3nThbTuogUT9GvRbPJaN7385LIZM+HSOSKTK3CD94Lpzq5Bj45o6Y5QC3i9av9S/
W9yS10xBVlB3wFojwr0IzMzUk83WDx351ShSpbkK31Yh2N4NlyVaz6ig8GIskX8zg23vR20zeCMb
9RuhX2EN+hlXlevwJXnlcw17q/NxlJZICSFVp7oT/Xz2Q+4LzLD5tfBOCegezZNHOVtp1txtpNvL
79cH/zpa+98pb5Cz+7qnNO8ecnaGLOda4LYb1q7DDstl9qpe2gq0cEfNZjKEmvHjndctIh/snnH6
AX+hWoND3Jump854LPcovA4FEtkVJyHF98k455aVZo8tcdPvjW9A1WnAr+GnsJANMkJPHPN1mDHB
Nul2vXh1UULDCydoS7AUTs/+h9WD9No8s9zfbQ8nDJeoG6S4ceVoOenUD0fe/tWp1BqWompDkz2/
6I460D3obcLCS+642mq6vH+7EsfyXy5/Pcg07QE/40aOfUMfRF2ujTpJ/alCPO3ZNRDl3tEI4Hsm
hTI28l3G88x/GY8RB4D4AwKOI3LBePsyXR13N7WNxO7xrrOKt6Csj4+GsAgulh3vItatMSDeilz0
CKEMnMRub/+hh+bAXrZfgzJZtRxrozIcKVr+DrK50z42sWmx97VLuHADif5aF/YkgwI6nEg8hkSs
a2w8a38z+/W7OqgRzp5NAgUSepbskFEmH5n84TJwp5mDqhs4L+v5wtc6TrFAxuxgYkwKSASOKwFP
/jojpWvqPQ5k0g7jeyu+dOGUUWLhtqGWv5JDpToSqfGyNStR/U/6yWp8TC88fXdnitqkiebBYytb
RLZGrRGvmTL4AewWbh8ygmtdLiGRZjzuh9kOZ8K4Cor8G0gagbXZzco8KMeRgHw4/Bw+67TxLlCG
PI+c5aWzcZgfpYvtnl5Ij4h/3FjYYk7uhzhYl2y1saYb3SYgVQSI9NPNbjO0rj4Muo3aUl8YV5NZ
hYnccTue9gKy6pgphs76eon1+hd6WdZHiarB9zo+8n3rwQ0Pb43oLqUi+oj7SNpTEzZuub+TMdLd
uEfzLVL4rv6fUZp7jFWCe2yFSXRdexE0J4WWCQFpCwQfcQxpQPTQ15tcpYtd/mYBXOK9aPA2tH9z
vbhINcOaDUFGF1u2oH+X8GSs8ckahJVdgOMhHM8y7kCb3nJybwLvC5P1eFjeKnQG1Ne+V2TjDIdE
COCf8rhYQ66VaYfFxyCAJZ8h6uxboV/ABdMW32BnaMtvhQD8+VN8lDSOQKLe1mvpGr8BS4Y42T5V
io8rhPAsEpDxwNOjgGbMzRtzFrlvYLy6cSbOWxsQveJz3OagIQGii4q9pdH25Wg9nPCZA+BIluBP
iStaToava/gYQ7RAfIk+1uZQ+Rl6hAF0Mb3NhDMJDYjI83iL4IMfPQSGrF8PZ0EkbD++mertGvbK
M3AmvcV4sYTQ7iQUlINWRmSCe5qgsjD2GEndfk67fUTUrSCiZEvEqZ5FidHSMd+U44wGzQl6hNjK
VJSAj0VN9GWg1ADLv4FrdiCJyEb+iCDHUpKRlK1kCBSKiSuXur6tomYtcbJHpk7Pp0VBBGN8lteB
CVrCkgAw0o3YzB85SSAQf+pzBkzI99wTYWkM2tBjiEHH9g+vuv/VawShcdkh38Cq+O6k/dv2N9u9
GT2mI+TCo3c6ysXrgMxvv1uvkHccJGDlI3IzQ/8s1S7b3YCb7c0G9IeQSuw1BMRlHTtVbx/s4UQ5
fkdHwf8HYSqHD1dOZpF1H89D1Izsm8XOtmKWHqrHgn1o78bd2MIQdeIgx0gPN9dW8M6wtVpSpYT9
fCagSYkiEtDgm6x2dpI0s04dhzKmNlt6fQmHtAMSyuEO/8IPlb6ZLePgQ3lvlh2pzGCbMk6I96MK
xJJECWV7RGTtXHUpWug/u5dPLq/3Vj4oDZWPjR+vmLTZtYxygryttQFDVKA4ONB/lAT0pNeUFjrk
HIDOeAsaaQdvm4zLsEt8oddfCX3zt1syjRNI6Fg8mSKmjCfn7VM9DiKZoRWdTLqpA4Q2Wk/PnUeO
QjVkZLrAPuciBC866AkDJNPhZ2dvhpeuUxaGAIAPf5rn0s8GWHo15aZvJN91Ip24pVRQ0i+ryCv0
QerWuI0Q3s2IorymDH6RThiXcRLslvJlYkQdG38QYHVscSl0cGD0bwljQDdrt//pMehuJ4xEvP8E
bVq6hDNKPgtScD4hwrF4FSnIi+yGIr5KweVANAnd9FT02URiWAcU4jb0+V9U8y02vdpltLFWCOdL
w5ESD9EjEF/akgFH5ehh3RweFeJ5sGusX2totQZzTA3N8PGHjvBNEZd+TmMdnp61fbKNR8gT7IvW
hdJUQK0pBjjTL+4xBuK0iCvOcHkc55iBG+xk1x33jqawvmerxd9gZQiHE63jcxKRbHTePFbREZHJ
+sLLxA5/5hqROGlvmyus++zgHCzg+q9kY+gh1zQcfX2gX6vnPgZoXd7U7OUu7sDgedIm2n3/KWas
pCX+f82MSmsbNGGwflTjnAjqQh1PWK8sLj2M/OkUgUNhaPWG6jFvnxiCZJ4GFLqHM6FYiQe3yFAj
NgWsyVaWKfN+lmDNtzShCls2tn8F21jVyt/kudubFekcWO/E+IRNhjX2AAzGV6McY0/EXd2LenLl
A+gLdGrbcB2Ay8pOK+A6Hmamk02cXcrOOqex6Loz6YTWTxi4pxWvCmxCAt1dYiHzqBQAAOmLmV3R
7PxJT/3XvWZFjsMpuoPpl2n8TYtzieyEeJ2rnQ0QUHQcTdqDtKJ5FxEk8lJmXZTnjaIHt+e/5j9P
VQ96oxzw+tl0UK0lHduN+DlMYLk8fw6UWOAWaarUgKLZapRhsD+C3Uzrf/9/3Cwmaoa5iot05aA8
o1M+oez0arrnMQk6zAr5+DireYu+z5xOI08w9J/9XalOdku9fEpQmmidwWytyVFIF+vWEF0rspnK
cP9Wufk8bwfegKDTIEjilxCNfBuAHpyMFxkSLWTueDDqWXeaH7CRBBRT+txS+F6P0SdGbckj3XQz
lPLg8aDq4AfECNmXjNyyb7aYkdnVGocMhSnw/287Vyy5/P1a7wA4+/WRzTNT1ykCE8rqFwUdIos0
UoOlncs4A41tBbcqLTxcqx0lxUl9afqGhAmmG+iHONZk5oLgWP+BGSivLONNahJx3hpI0kcGLc9p
W8a1ChfMzJIxIx5U63sH3fY0Z3vV9RPOiBw59XEgV/Zhfqb614fGddZWiaR5gjAdC0zMzSdeCgeJ
yjl1fIuits3EZCMROBpf5rdwk4Bw8Eg6M1HxKucLRra8Bmw0CV4MxjV/HuFAgQsbemzTuHG+EbSn
eAj4U5xg0dNghG0LN1IoKLXO91SqZe7yRfq/+i1x1EafTl4+FZIcI6spkq005C0Lxqey9d6zZpef
ZtU0n7ayyt9k7LXCIY+Z058+MG/ffLR0tWy9TcTOn4jNfUM25uBmngJqkT8KuN13YyiyxbEiQbN1
LaQrKRJSSqZklmbNf54b3c90k1C3h1W5iyfcjL3RqUlUkDYPIdyUVSLhL/TAn9MQ++kJz4mpRn/h
Ee/+JXnAheTLSoMBSH3PASahg+7cqwMtUecVwnXfjSLqrgZxkb3wFSEWcYuO11LIecuY43jIKjvO
kZiCFOlpcDwe1+pKyYGP1dvfQSK14brKNTS5qbo1pxTI5dDUWnsHxQBR2469ORuYnDeVQehrNSq+
Mu1T9ZCpx+mBx9CIkGv6CEXl4uamnwRDMemIUVFcY+tF187vVItUC5zS4jaN0L0OqzCgMi94D9rF
utOPQyxM/a9LjPfJGx0JtXAG9FDG8lRuRfQm7P7fqFKBCo5sPbvTKfpCpyPa1xG+e3gSa5RVFUck
wRm2gxfQwQ9FTks3DWvaF1ej/zni0f0ZZFmqirdFuqnkOIgnU7zF0J5Ztwot+0heh7KUSuAKvWzG
Fyo6HFLMPDPRqowVhhSY4vBIdwOxSauV0MsAYVV21alh84HIq7Q3pkBN/zAkKUQmltHNXYjtbmrm
uC+DBsIf9zN1M5vK6c9lNaH0SnYjMM0Xrre0LOfNXWg2J5FSsPNCaVDklTmjBiqoYTlOKnTgy+Pb
A8csu7Yt5LA3uCdznoz2gmCH4jh4NZUmSViIEHMmFSRqEIUrI/lXU+5OMheEerKID1R2Jg1AlBMx
VmBCZYOQ6AL9FdIMdI6j4D/5Fqz9UM0MR6UQH1tIzgCoVChDczESeGoJESekb/6TWUUPzB0EgCBB
mpT3ZR/kvDFvTufM9jmG/YZhUbgPwyhxcpy1vb47Vx0gK0XtnP0k4FM5VMYczXkd4FJELQT178l6
tr71jd2rBQVfw8gs2mSWzoenIuj26nB4DNiTwbXCXDEUiOsTAj2+Li7M2ZN1eEOJ28t3BXoAqfEI
rzifUyysjPiG4PVvqfH11k5ub7zLJWRBF7VBr16u9FKR+xjG37LoM+lW9xjMGYn6hhX/etmQqNhj
SWqfUYwd+Lz4E2HkIc9HznDJzFxRTaU1dOfnw/9+Nh+Qtr5ZH8CQxYmUmit8lHqrC+ZaIfuDlpPU
Hv1FIPgu6S5saPUt+ASOnFZLcnIuMqG4or7nfnHF1YUnl6dpkqMV1N+8kjXo57RCVmqMzyMao+GC
vdocQAd/JIxihPgsUFXjWhfwdJ2gAsJ+e/f+hgf32NvynLA3vdjSSkUpg7ea9zmwCJWM/OYEGwQB
lNwVs75AGvAOd0QGOMWrpYXxgl+itJ5QpHNYxVmXWEIUT/rjECVinjWP0txC8L/119pFD9bBoYTT
kEblfY/rz5b9xG9FP19o+8USZ1H/Y78H3h+cWpp6amdj/1NpnpNcqfCyWEQT5qtbhvUXB3QfysKz
NPq4PKGIhYwFcmNlGpE8CC8lYqltVGSOXb9aE5lyP9NC+iM9DdYbBMZ4/9H2JmevO0TQHh7xL9h1
1N2RZQgNAZRDmlyqB44Y7BryEP0a02dmiFKB/om5g0xDNyhEk3JOuTVyJFm5GyxukxSXqPGJm1Bm
SItuuom31vJxJ+dl0H7XPHBAp5B+V1g6v+qAEJxwrjmf+8VseeL1QlcKCL18xEYhZe6hs7xboi6J
F9mZDtJLcVT0yFcnAkrxfDpH7mSrH9fv+7DOQWjUzWl0dXxdPMiTUb2efbHUq1XXWplJJJKHVGLx
R88w0VR9MZcuFALJJhZnBdPoI6iAvqZEGzH2NFMFfD+801btLFWtuyqD4GOjDDPf46YTcWFYWDze
Y5cmRDxVO8WCT5Y2+IeaWm6i0Z6vyVpp0tyH18gfqdYRCjuMMbVJjJmd5BIbt2ynhYdXTTy/pkt5
1H4ywDl2TLw++2GhRIE495PJTaDb/pPQn0Dl95DeqML9gPV+A8nIxMwAI3l8ZmByUfAaMngkGx9X
zIAf6+t/J0vvE2xUpGizrtw1rqzt/Il9FCFXNyRauw6gasF5y7qT7zcNlmol77fBnWCznUCtFOvV
QbepapWXXrdSe9/KMy7Hzw2MG9UsxzJlJM4Unc2xykJnxHZDYF+oz7O2ji5Xf0wrWitag+la/qeh
OhngCAKKYzsVJ+QvczAcvjRN+jVCh9J0yYEurPbyopFM2oBlSvVVEJTQBRdjxmBG1zPTGxIQEtVF
HQnphCZRwVjmRTA9Y69lrZ243+5GnHnp9GL603iw0aKQI5f1NjJez/tZArWqNdB4dwhbOY1UtwT3
MJKiLetHnFD0TLfW3t7Qvj/dZgqoo86xbJnLAQJ+nbyL+8ujqLn4ex2+vplhFJuyEzQ2JExGJSLg
CvmXQerBkxDo6L1QJQkBV73nAv6iDtC28QRIwNWOa8EB8rc1cvdUYPulaga704wAzoMCJd6BcQeI
MHz7HYRQ15wVdX1JLDQDhUMFtlfurp8NX7g9ZiVrnP6s3i3i7p4AKp3PoVNwsw/RjO56lehTW8S1
ho05btAfWAtFTKeDPeu4ZmwvdTND9M+J1TBA5nfebX1NpLHxfIYOGLrR7wZdb8lM3BoJYqlz6Wao
OstYawtgbd34nsyz6rJl74FOG0Kg7CDWYt0/Vii9DQiw4LD4GVygev3NrTl/G7yMuOb5VYMbMZMM
yOi7RnTKyl8I16tes4VBPuws77oQ+tpiw9xZDv3Qd8+CO9Gl27Vlq86S/7e8Y6qkV7d3CrKbu/jm
orObh9IhHRBcQI1ayxLHdoF3+zkohO0WkBe0gpUdrisjc+iPsyMBN8DZd6HQr4wBOafHQn2AlqYy
XYXbvFL94Scj6FxlvXKJKF2EGTKDJF/G8ifDwmWk3GTVsvEvmo5TnCAupFlIfvPhf2oGtwJaeC77
xqFxORb+xPEC+2iNtRv4XlZzj/qeavswezO786nyOt543prtqR8BxfYuZPE/7BVRIH4BLU+9P/W6
P7EquqgykmpB2BzcI4aiC7Mo2jb9/dslW46ardfn1R5ZLsUunSDAtbxzZm0HYi1/3LKxDVzI8e/O
OlEiffWUFXCRlCHn2AFhC2kS77l7K7GcVn0Ia639GMdmruA9JDfry7qQi8R9mDx+SOdyqOjt2I70
B/38MM1N76Bh04aLhot7DfogFh7iCxsXIM0cuKOxdHMv1V9PFm7ldbhIoweoLsH/vFxVgIVtbTPp
XNbJ23e4S9ZI7tY9vCKlbCASelYHkL2Akn1Rfhr8/Ev+4n/sFn0yGbyx3vZybG3m8RinzAzznpgO
Bl+5Z0tZWWHgrmVc7GaSZvBgz7z6ScW9sNjyRurW16cxycZQ3W275W0t19nzKTAuvAzhce6RZNyE
7c1NFyNkstUVZFk8j9FMiJM6qBQGKD7JLnY0RNjct7AxQEJ1GqehgekmN9Sp8hYwdjp19ORUwczM
fw3wZhSR/S9CWYU1xt3n9TtapXYo8+Fg2leSn/Y/LNvBqEw32rJrFf2UohyQi4EKhiOjdokJp+0c
R5461xR5ojcL0wcW6+qqooN/g48LDKeE8nxxDPFQP+zUM2wxPZh+qFqCTth0Q8RoPnHP58PM3d5M
cXHvLKcEj59eAIElqCoZQqFHI3JZcCTeCQu+QdG5QXRbuv/qDVDhUyBhb8FTw3O9NRFp78+5qCfd
7WACw01bNETp7bxaqx2VTphEe8NRWWH3QsNGok4ei7Eql+G9Eka719GiUX8YtPrd+ccB/Z6nxsLo
HafGwyJLJi7CnLqUoSOkkfJwbLOxD3zziMmEMCsepO04PNC2kWo34Q0YenpCNlQjE1W8Im/+jyud
L8UFvWOddxagQZNST7yLeKQ4dflIHCbc+A7NNMrD0OlYJQ3Cvp6bhFXwuAeIp1fRiS6bOovBX1EF
NctTtiRI+RhjfHPoxaTOD+d20F6+9Vdkuwtm8c5dCgeUc5f8DHa0w0lvd8H3kTtwfdJlv6LBPAfm
rJ5yNbdty2R0DS6Cg/W2s7NysfEhuMzaoFNg/TWW3rXdRQ7hY6HZnDQGIvdqqvNyEA6XoEnI3hE0
FqHgXpoOSNo8E/xNQ2YlvArtqMtNnKINfkDNSrGtERZsJu34oYkLgLqk5K8SNSNCU7uNb//gY3QE
63gvw9ItCg3sSZOeuFyH59RQxD+W4mv6rjZNeeI2yW4fYuF+F7Dyad0DRWX+4GZ8+cnh6dKnJTBy
K9LuP4JuL2R+znKD9raTIcvEtrmKoHEQIO7NAM2PQxfkWi0nf8UcgzZ2VRi4guQ2SAq5bUsYz5aK
HI4fOGxF06ElxqXsGwQH46Mq/P7q9/VzsU3q7hlpphEHBnawbUSf+CWkeB1N/ZqtwvXqsYkNvz7U
Cs0TMIIMKgU9eNtqBnZSdA/3PYTVs0aCaRh01mcLBbE0p4BzAmvkXz41IaA85sKoD0xcWEkV1LNe
3a6hSb2l+yAkrJ06J7LJQ0sBpybPTw3qmZBols0njMSwQ0LYlEV0JPconfzM67uAD9fB14pBp3PQ
ztqWmQ3GMNUSZZtKt7Ui3PKQfoFe50jKqBxaec8ysAhSc0UMbOypCyQNTEwrAzLWje+3UgDvi8wB
tJQRC6so5euLU3Y+j1XO07hM5T/Aa1cd7m/ExPmr2GdB/u4zzfg2jkzyWNSRZ1VvH8uuU9un9yoc
HpWJahuCT54W4J3oVAbBNj+awhkWStyAkB0dJRiAkA+f1YDWR1tG1JMx0LeR18zsfnxolq8WFwUz
Hc+DY90nI8PZFUbaDHFv20Y8wvPS9/Ivp9EwyqwpQAWN0rEAtbC/q/xa3DF3DVTrEHSmBYSh9+zu
hHeNYRSA9yBm2aFIdpvWCiaJF9wqMFMPg6R93dsOJq16ufIgUOdMGw3daLwVsNhU0LjCrgiO0XL1
ywdIIPByDHdPM/x2B1IYuEssYKYwk7Q4ytjUU8Nhm08sJ1wKmSwe/sssWXQR273/PQvePDd8a8Ip
DFvktVOT92jLfXV5zufze/eMaKiW9vPMJTc3L6oppm/7oafREXAedWPm9gAcfYl1BCVGN+bEkQ+P
utoHKJUtcsmaNGYCMylFyud46usPjl2L3C5JUpntjh78VThMHsxuAWFZXCuKHo/K0pZD0+00meCk
RAELMXXmLNQVlzlsmQx8hdc8FiVlftb0GezSTFX//DNtmi0SecXbT1I3AFEaRuX5fmAAFHvUfYJg
2q/s6lARIBHZZtd7CIsTnuyGlu22lqkXBj42I6HI/d5HBxVSL8ERvM25Wwk5xrWzlq7euCbyFVfX
ZwvtbkRBab87+io4leEgu6EthbKeyUim1BEh+ADezU1VpB6uzRufvhc9hzIA1CpO9rOTQ++Eq2FK
4K+Ij2CHsIdy8B7XR3xXHlY/BzRGAo8GvCUQQJ9UV1v98m1qFsMVZAdUa+YMGunNuBGX3zT98CIB
pHZax9NC8aUNIfuNSVqvgS+HoAMstiBHq9YxSgc3MzdeU2lIOHkneO4rXW82/SxLPLHqj4UjgnrO
4dCGzRzAkl4T6TodGt4eGLRr36Z6WmU7w3USWybUktRSsGq0ACU92kIV9Pn8oezc29j9OcKHK49t
PL/WHBxjiYBizVbctBgSJChMuNnGCKbS102/W1rfCeWrbM3R3GlRgF/o08pXHmmTAqMeNIeC/a1Y
CbDQjVztJRMeD/Hfr8GZQ31FINXYhoxp55Lhr/RyouRoXAQCaVlJjD2kf9BRpXW5uBGFH6K0r6r7
EVaxhCyC90N2DALhpO81YrK4nX/4sXNJ68V+VrjBFQIRa9I01NRsOgxF3E571w7uZtE6ifGk4O8q
kPGO2xD5SxkSE6KTf30oVNboNDByOLhAJ8qVoeudbgfeOjxbkaT+2nyYsi304c14FbmvK7fjBkdV
hF67+BoT64NI8VG9E0ss5/hWuj8Hz437BXEncBufNHyQgWslmx+s0LuFgQ5GaXj7+5pQJ7Y02NWb
4OQU4bxIVntyEdAEKbZ41g3xuiak2wm5wqwvNd1HaugRYQsfaaCqQkLPKPmLtsAHBCZwxeq67lPt
wZ/90ICQcafgXDdQUqjj4my9U811zYdFqRh/MdVBPD0HgmtihaqljaJRW8w6cNC0/UEU1w667YAu
d7vNYJDm1xPDDiABbk7fBO2y/G0gsS2Xnpm/zIFCM5sOf+3DqZvQ50KFZthlIhbwl05M/Nvz2bFL
50PCRog99xYIl2sLLno1pKyq4HkmIhKKp3lkVlRF3Az78jl9iWjKNJDhXuPF1Y+liwlw15wAG7jm
aHfNmt+SXn6H4TGTwVANocQdn+vnaKQFcBQFZX0ZbDE48rgKqekeVUYAOo5kfKiGayDVffkuAQNL
yWPNf/qMSmlzfjPw3gPoBrtqTe7Fm7tqfd9L8nlR+0hpQdcrPyQlnhujF7pMoRF3Ov9uYkvJUOQS
+MsV3+wAgaDGW5o2f8+DiHa1L6WjpWu0YYaxbVxH0hSxbEd89gT8cp1SVuHgk5d2CpybTfg9gETP
0lNmcCwymTaHW8eSxOAdu8Hfbe5kG0lgDo/chzI6SmScHevUGBGVc5ZwkafcEfwD+9busIs81pgX
+Vz6S/OI0BvlkMPv/w5+Ag468U+DiDJkaReFP9lkSANqqtLprLRCv/9/zsJCl4UxuyJA0bX1FJuk
dDxHRzIH2bnGTfXnMOMTrlUT1WsJlWcj6KOIvoq+ppMkD92OoJsbSy96xpRVNe7tA2MUPMAAuFJV
IgI7jQc250WIQwLJxBGPf6auhPPgr1t9Z43Rh+oTvvlCtzsYQdSTfvDUyUVThAS3M6QrpbFUAPMJ
/cWfVlaBEpttvC05tys/b9cPfk9zfFaOSnpkE4B/Mrgzg/HFNV3Y1odWjG8nrTrIfBfM76XgosTy
CfUQFCkJ1Z4jhJNZxF61VmwU78815mb/j6lvJ1DBp+SmkMwk06XhLJEa7ypxCaviKOLuL0iuSH9/
sboxeuS04W3Wlk9wBTDqEnL0DyjSceDaPTouesiRFqhg24hyqFrTmlWnkKXzCFoNkMrnFAdWvSE+
MWlhaFpYQWRoeuQ74bB9XpkFkLdrq+IiZtHvLxoBY6URL1Ea7CuBw/merlM8kTvw4xsym0uvCKjE
+C3AeYPh2ZKyFF5X8A2E6luuSrqDcgnYNg+2jUJCkhH2kKtz6Y8QHlbBklEynrKFjrUehNpr2NRJ
CRrzsfbrDIuM4WdAz7baXbIVWL9V0XPdGoGlBRWZh1xtjnn46Bm4nGnbocQLSm5miLVNtv+UNROm
pAZaAzG0e4W1BKcaasBwsTXacojVLDLtU+yJSagzHSncPcAHiT0YMBh4yImZ4PLq/dJMHxoIzIvw
NRSboR6FivD8PPRm5VizagylyLj8fXJ/4o76uI0A0xXcs5YKTVfI/f5ptmTLIr+8Wkb0pPIV7/gP
aZME5USt5tlQcnTLH4wSdwUKOMJ/kuaKLB2s6zTvy6mA4S9pE8aMcvvmYHTXY5erwhDgYfpsLbWp
DPbMlc5HUZCjT8fmxD21Aasf4xwuz1E1gxcvlWoDxVQEZwPgVQk134dC19/ZqrL8sZo7XStED+5I
X0kqLnrIYeaDOT2UuXJQ7qE7HrfUDat4bXQfMr3C6NZjIFuDs/HMKY2wCev7LM8Y+nQ+VfcneW6S
uvfNXWn9M+pnVD93h+SXURwRFKjcLbDpVNqmxEqLCtRuxxqOHdkEskZMA0MS2dZu5ngvJzLqLZT1
/t+Jl4Jtx+/8gCoXxB7RnCJ696R9gSREuTTiW0ZWvQw7Mld71+7qD4xQEcOt44nzC9+BcwP+gtQh
FfaMjmF/H8P73z+hXEjRHL0yCD5LDxWJ6aHY7E6XdQOl//zejuytlS103TMhbyQqk0lhxS02/guz
MPucfI43rojFlylkmYi1ZCn1eb4GqxEsLu6KmEO8iOEkDDYo8V86fWRAG7zOBi1EObO9ECL7oSBK
MpzpLMPWV+bPUyNYWWSR6/FiXl4WPBAFAW2CHkQS1KtaQGqIUrCxOgwhiS0LoBxXkZn+xP3TFnA/
8ZxJjnPfTlN6dbmdmaQevjcgignjsfKI5i9szG80RHOmEfudDgP3QsJ2ydo2bAGzp60nb0D7OmIm
7pP64qGleNmDem2s8/mP/NZlZvriZoiJkwu2VHYA1+N6m89rK3nDThhwuFa3LBY53E10r3nU1MU7
lotnai7vGQ/tBtjnR37F/W9IB1XxzzeMlQFuxY+vtFtU1C4uLiK/RpKPzdLT2ALts4wIJzsi/mpN
gHHU9gjgYLnvr75UKatVJas2jeGk7HE6oHwbTyFHTcFVAExHyo11Rmu4WW0vVYcC5I14tfSVzut5
NzwbKJ9891OTmGRBKpJuqWKlvT6SMOWOBRTzAfliEZHWE9WbKNNN+NEfMNYZeUYhmn993UgACIHq
aX5bZZvVuIUFbX8RbV5vyq2QKgrh4SwFdQNbiGY+VaNRCchYbB4KCLWSylPLlLrYDVIlwjIMP7jt
ayxSSi3J7YSnhso51NK4ok8MbvsGJgT9C9F2+hzLEzD1h2hZFJNKL27HJqLOUUk3Ll+2LaftUbfW
DiEzar3v1WMi2lYXeLL/j5jp7A8hourZ51IaBgZzm3ODEfJzX6/3x5pM31y2MBzLy9pAKeHvCyQu
qqJpjSL6eubzOh16mKPp1saAOh14ylW15RjOOdTYlQeamyRtQV7oKzl03RmUmLgifQAglb5/VyTt
98EH5nP+CuMUSSwGwOGYZDu2QrFrcZudWhmHF9pKWbO7/7yBH5JfOmS6KBtQNR7g8sigRRiab8+i
mxHpt4GFof480yvqiBi4ttRd2337SdbChsv39f0USvANyOHjby2ZtmzeH93xkLlPbXqZG+ID5eZL
GX0/8JFq6ZfzaJpecozoW2jrtMAJMaVKVvbKiQjrHH/7ddRD3W7065qmYDV4ai2ktjUMUR53Hg1W
cChynoAaXvAYfaRtY9UIWY1W7CkOV+6g5YnGR2t6kWNqCO5ST2SYnnM0EObdYSHJrdT7Y0JrLiDp
Q2TC4betTl6L4eiWv4iuA9SAaX7KdcRl6VKtdeI2iCLN1grZ17qiVRSiW382jm3gIIv4NLuF0Rnt
h6jPL0FRiJibOdRei+tj8MrzRI/aifyRKItoIIFf6dljJAfmH8he2sqRP7Tyk4Wwpg+h89mGA23P
I7LcWV5JyUaxtwwUFFzfDB/1QYnz90LFVsN/xH/2jkTuuXy60lHTjiGV8uuXjEeoQpGaJDZXnfYJ
9QfAAEhalfqAwJeLFgTfyl7dObHFf4qFgQ20S7NfqHW12L1ERnDPNdz9ow5Nh1t/Wm3FD3WAyspR
X3R0suw/td+htexrqV4/OFUwA/11HlLkpmnnp3wqL0PxW9scIDbhQk2hYX9ElCROMf7KW5zbnmRF
L6nqUQ1hUeXfvZ9HO59vQASncjNhi6Y+1Jyidy0W0DQv0ucqlzab3YsEqYXx4pCaRhqYSdXUldV3
8JoTy8QHIOqjiRVHDNH+zTA/rVUnL+c01iYlpUsA2lbDlqXd7T9k/eWmuzbx70JlDBotEz5T1sJM
454VBJtC20sq8tEg3BDGQ2RIVDqEeE5Y0xzTax+q5503x67jLyrp6avv07eGSH+bqcB3HOrurtnr
IDt84APw4dRp7100PcjxrUgov4Yd2zKbGC5CRVyFbyOt9kbKAC31f0vBugcLZyS4g7mEgGiBZD2u
00FsNc7dPNIZ6KXCwKbPp955UQvmWrbLPXy95KSHHVq59gh5ezzPk4xN0lb4Ml41UNzwSq+iAFMj
O2myS+pr1N8YNtQnAO0eq4wBPk9vYRAKKS5CMxG3wFNP3WO9jyXxfs9fopK75dfHmYLUE1EjLa02
Tr797JB7E6TtXnXVMpkD/QkCA9JXM8RSYnX6NHsKFkH2j24dZkWhnUMPWU4ygGr5fmYQsTw0BvPg
g8BFXlTggnMC9SQhg87mbajQT6Xlon+bdpj+bDXeEz7exv1AVz0JaC3YRTE6LlGCeckDW3Wrgh0x
HYu876FqnANduIQD8XaG0bKzA5320CH4LTSaNyZXFAA2eDazBwJtQwrAIcga2QFCjPQDstBdAXgd
F4FdO6Vrsi0eONlYMmDl5WmB3ZUbyjWZx+L2zCvBtolLEH/hINeR2XeQ+VC8Aa5laggq/HLci4JD
GeqL6PRAuGyDvJyWTIlFW7g8HqsoNvC5zdcfc2AEbuXNgW3ZZh1Xg3B+9HpEcYjTfoW8+Bxu9XyU
yUK1aRmNMDQ9NCE956S6dSukcokBrKjPacFD7bYVUxIt6Nft+vKYH8tQJiaxVPMZh4E/G/euaq5y
KRIxPzepKa6xHQHQMZtHOz+YGAlkcUVJnJcFoerHByNa6NcL4C4/TdREqRT/Ypqq4qkwhOSGdZQR
EK58g0cWRCrACNjQEtNIfJfYZUW3R7RM9681fYtSG5dmPFDYsz6TkDeZqGRahz6X4gwC5A/XeROB
gUnZKqF42F+BXXspj4Nh86V8x5OSDLfG41GAihfZNeqeDeaCT6bfbtPjrwMgeeCtILof4E+Cfxcr
N5BuUEMiUkCLOtrELxgAsXxZdZc5NW+Dx7RMkLc8KczuUN/tEZFJ4KuTaQxey8zCZRcXSmwzX1AV
uWK0AkfIV/DBJwksfHF7i6ek4gPSOxPg/knuTaKyg0rjF9LwxlSJ9Y0MUEDWHE0E1cAe2noL55RB
qKj9u8g7I2cl0U1TBw4J1xQnFaHtEegjQeXh2PqbmKEhqQkkz9jvsJqYIDJC+NRJS/vsxPHNTL6Y
eBEImfepmMwi+kqjG+IryonIY+84zf8Mkzm2cLzPt4PaLXToquD1/4HEH8u6bwXtN3Di8RldvvIc
oi0cccv2VIAG+fosU2Sj8RvffORVE3JHWb4HnqvXQZsN1s3K3ykDMfeU5b/76BabZHqrrO86Gnv0
Pug+/7RjlbtXjXYk63peoSIOSf1O2bmKkGMrs7xNeqmZUWBKgr1Lwc2B56c9Kny8rGKkgcV8/P/y
CiHOgGFuBhmqrE0/KglOvR2pvttTCrAQB0N4PpqtYx5w/Dnjhtjmx6z9Phs7Nx3aKE7uEJ6T7RMY
xMeWF60GprwcNDuBm65D+YXelAx9ntAUCU37qhob4CwqdKXJ2uAol9EyMh8oDk9uh3qoB3T9a2Ng
UwuOfVdJIZn8FaO/QmW17qcaLqstHN/j+2Vk7Vtf58Jl67o77Qc98eGXJAM5LEVjCSNHu9t1rgPK
CUB9KTetKUMMwMzLjMlIMsOPlDvMkUXV9Or+Er2//SX8uZDWrGqwhCGGMY4Lc07NGHECCtfkSj00
a2nLUxWQsuKJl8ktKttpHWL+e8Rh0XSvzUK6wz1vGb2Hw5Kat9Mgyyb0MaRExV6U2TxCe6pekvAC
KRs6q4S8FZPZ7iD0mLqCzphYU0bbVb3mqZPbN2YvKtQ9mmz5S7h4XXOJvbO55P67Zel/slY0cvJc
aGFNVNT0+b05VW9enMpn9GpsMajNB55w2IdsivPBBUBwQa1FxLDQJVslDUngJVuKfvEMj0JG5K93
0KJgGhLpsu/sQNKuj07tCgws8N+3/tMaUTB8NHt5sJpt7F7s0iwvtJTA8r5gmjWS4KnYlMEFLzaJ
dNexsKMXQAW1cSTtkFDX+aWC7NhTc/KbScCc3pNhM7uXECdxq3JvZ6GVT9txyKWRWDC2B9lBgX+n
qMAjQXt04zIoAcyIYBSK5487hN4xfSjaWIu/wq2EsuXRvaI/tGCOWf+qsRCDPOdgNbG/s9htnsXY
JpeWZW5Rpi0rPOvTUAUKSXJ/t7do/Z0/FMA49bBjWBSXStUuq/v5i9xIqOmtsAewSwTvtTJNsHpk
sqXbVKaLioW7z0lY5DFs9Vg+sEX/kDczXZtCD7CWs3NiNxTUwV0+vdclhFxiU9oJYIH/mDi3SC37
htUi7l3VKY8vsqJIP/gjjsFOMmLzINkh8wmN0E81M55iF5mZIvDP0zMBoGwOUlbwNr+EdTdxM3/r
xlbu8pN/WJzYydrk6vNge3kvALJ8BFQ1nNuQzdNe+JnmfAExyUqFnMASKd3/g/dXUCURhg8oYxUk
1G4e0vkVYlhUTNPqFuW6c7p6u79iKApmwaGuE2lEepzN/7J3u8pUJ/lC17j1qw26tHrZkbEEP5J/
mJPSeQ3DKVqqyPraJKEg/2cQTHTR6zuiFQoEqEFe7gdjErFk5ArHYIbSn5l4DIn1KTFY8Lz8MSvk
QWFHOHzhRbvUXChWXMwZDvfzD3vpdC7hkPqH6YWCwgDEv2SjMnblzrv2gZpIkEWeAKSbBfAY40r+
dtkrz1A+l0t1lT3XrCyc2xphCBzE1XUaaYPt4OUJ9Vzor7Y8JTMImQ/NyJjcfR9FHpVch0IkEinn
ger70qRazY6V5/Sjj2VH0swkeO5g1OacCGtkAR3f2Ar4uREL3nidaoPopbSmqa9LjvCWHraHN+bF
QEzLAUYEyrTQVZCR35I7x56RbrrSL16ncepsGQ0ip3Tc6ibU5ludR+xJE6wzKTVUpd2+1eA6EhEm
N8Hcad3Xi2K0/AuiIMABXi9fa6F8fOehP/EJpaZ68WWemWzHj+hVBrgjVOy7cnM3pDrkI7A6txgM
rgTU3isqfexK4Jb6GoLxJ21ZrOyCwVuIVZNo/IVRPRjxLKcohwelaz98D6C2VnKleDaM//LtLfjY
mZvc3PHHQPQBT+PezeDwpisW+uDaNuoEt/jDZKXgwTtK90oknGa3zXlSbxA2d4h9kWSvo4qey2ps
zC9xWJYzcL02DDdYQ0fIFZveT4xdzTCFTZcdFige07vcl4I1Qa5fI0zthXWveS1CKm/DZpi5qNd0
MIADldwHFhvnirUAFiO082bgzZbJZI2x9AhB9oGsSSCn8dE3h44YEsXK+ANV8AfkW9AwdJHaXnrd
W2wJLA6TJUDi9FEZsuOOBuPqkxjqoxVeOWc8s9JZ8rn1Ht76Qa7/9okPtbEKPbFoL2YYavZSQx6u
0veklPFy3UezM+dATR/Ul9RBPhoKhQMgxAC5kCTgGR6FD50twZN59U6ojmHRALLtqBS8LzGWBhIC
Gc5OSNgDVPV52LT122A4aX6y6MFc44/zIFhi09Q3cQe1FjhTaAE4uUG58Nl36dS7+tY8/uY5fLPC
NRo7ZjyRNw+sS1C1lFMjVUyyMrlhMI0C1I9RwdYMA13OT0dHFfahzQ+1ipXnQUkcthEo5ZUZrndr
K67KQGzEAsIauDhUw9LFOOf0MU987cdRmVybPApRSZbumjt7BZRuo5ENc2wPFLUX0PKmgLbqPTj0
xnscii2ayDvYXOi3JSFPDwP+fjSgRAz/lR1LiW7qm/mLTN42SKwbM2UVidZ2xS/qdeyTRpCLSsn9
WeDNuml7uxz1FU1AyxYOLCuJSpmnfilGOOnR83rFB1hzFtCEjrVDsUe3qfcS372ZPsqrWJoeVZBp
Bb7abNgq2VzxACxGBwmt/BXAnRMPDuUVrZqLXLnkktyBcVEaf4oatS6JpiCyuJwFfZUJnP/sgVHL
xJAHqHv34F4W1YnnBUiYXJ5GfIB+zrPH+aXT3pSDjJfaqvx48WEWmBCiiOU8KTmqPPPPT9TB0eyh
WILz/rfJ/W6fWiNp+AncurpIqEu97r8vTY4zjX/Y+g7TNMqhh7v8gdIHZaSDz+DSZBUjpSWo7+3+
SD97PudzC0EhcNGEaVxyRvP5ahlNa5g8dGaizoHpqn1n9seNWDDxKlDNG1QA0pbnFNOPzkzhVpir
0gUFI2MJnGnUlGkvn632Osin6MC4qulyd9St4MFzM88Jf3i2MXOePTN+tq03I4ZSqBi9vh4mdG3y
2YOV1f1YSHbE/0btWDaRCknGm9ZoTzhYxMk72LzEUP4/jEOriKYdnwYrBoAon6A3tTi5bGHhdENU
xovpn/7qJu8yrko7MsvM8bCHFJGia86dUr2Wd7PFQpLnW20ilDkGseOuro2jZ1K5alElRnCUeuJS
gMrdEnSMBoo0PyRA9JKlriOlVhJqoIB7TxjGaPFF/HoylQn5RWou1y1LvC71EMrfHEs24PXJfJiK
v+BFs7rQE8k3APr97Lbgu4GhRuYKssqhhoZc2+wmuyYfSWUW13Q9aRZ72MF3E4SQCaiK3vpjR2ZZ
G3g8BCw7QM1j6P0PO4nA77GyH1EA96mqEwChq+DZt+mKy2CQ8Rrk5J3F7WApgpUpPxadUom7xFrz
vX6wYveWEHU0NB2hzCFHTZHWlw46IQVLABiLMH5/9VKlczSqv3tb9+QSlYRzTgZ6bCdh56G2r5Af
iGUHueS47qmepja9RUsGN2U/SzBSMEAihpDiRUZCR7Rr/PQeWwI4zb9xGXxlTjT/Xo8LOVdqySwz
JkUdxPXHAFYUzNbFoG2t0Hbxo7KgBCEFgPpr7JUFUmas/NAAdaIg0T/K6UUyDjY0ztV5VBI+P71u
pV4+aB0pljg6db7HrvwzKmAj3IAw4gT/1VeubXuulKvm6MXYD814stmbIzWG7pVbPZ6L346UAbfx
WCsSVfwAcyoO6rQwFn+Lpeq2GmyuIUb4D7R6TVhFRzHlnCcGVu4kZ3nKWFjEyIzpzcTnqmi2BIbf
JSm7p05AyUo2oBz97YJkDCWyDuRK/Ir/jXy27PVM/dYzn3XgQPwjyYP09c1DNGJQdcSKlJeFqq39
shpJ7wqwmppHuQKFcYGFtJUrKSx2XqPdOekTxuSs9tVX2lgfOXcbYl+LLYa3yW3h/ZuDLZIPQRXt
J9KOTnB4MsgsCe331VjZ1VZMTbvhsupA4sNuo8c3CAutKeBpV0wos9DnKVD3TSgCccrhd+KaYEFR
wrg0RCbUNmSOpaXlx0zEIIJyslkGKzYfLckh2mDif/KfSVNzufXwvUesRIEnl0RrrK0zNFNQR2c8
frFwmcYxvdAyPQR9/UjDbCwivSUN6u8RsNImEu1cEq8h2+JwPklv6uV/isaeguRM/Zx3fapAquzk
YTtb7jfUs3EyD9TeiPB8UYPQ2OiTb7j6CYWYNA7IGxqKrRVkrcfUbPlnhFGuVELJI+48yLZcGB1o
4TaZXPYvsXn84t04pPA4bq36IRrO8Lmn+9TiAxr3zDQEAGZVMC2MkTRd8NBVbb0g8dqeVauJNt63
IHVb7pOSaW+6NOOY0L1ZLCSDBDDwMCvb2N4FbbUVfW8mtPoRARSJ0AKae9bxIMxWOGxpLKHRz6CJ
kf3RJFPxC/h03UxKPCzLxDOqmimHtyePrgaSaXqjXx4mKyyhgqd3sM8flFB7v0fXMtdqnmWS5IOD
lEs1KxA6AFFlGr89+6BywSurWkgoT9UdHSgwYaAFy5ruEf+PZv1qFKxgNVv8Z3SxsgW+tCaCktfi
obeVCZPqvprgj0oV75Sjy0hSiK49nJi/VByM1skwBlbtzioqPhLT4kVwqgLmia3GeEj356Wb4dEv
981E/IWjuHYpk9kZsDi3X7o+lQJ/QqyyQ4NmoKnajkKzuntZkAuHIO04QM3G7A53NP22OIcer/oW
tShs9HUADgFTYCxQSM28LYC4y6bDC4TAfcHuWx6TaM1QOVgDLAnxTcFCWS85w5hQwQDkPX5LZv0d
LWAnTMwW/LTccjiTXhxXyWrtqOQLJQ0e3ybwcOWxg3dRnHRgN/IuF2pgENV1YEe0hom2YgAInTLj
ev1WVgkrmtctBJaFsSUIOnbuaJC8oSsIXfUSMF67hgt8H4G0e2uOHi//pnmAfavVNAVve005++lF
kJ1XFJqYRZgEqfC4rls+3R/yBkF4FqInZ4whEJ1YK1dq0NmSS/y8RyPUBrM5m9b41mZ8newAt2Fx
9z/1QG0o4kLjWFhfanVdguZ3m1Sssrniqdbs09p9vuLo1fWFKoLcQfWK5s9G9RoPnGAZWsyz5ICb
k/DM8xLJsttTG6ld+STEFKARkHY1rK/9Snp/dUJVISfysfbIb6oM6b52QJhFR5P+BlcQEnbQdlyG
K7fHm95uLuSE1qEis7WQeOujfpt3Ifm97+6127fkP1APbSkO4H78Q8s2lFG5nKhXmHg23i0lSfhe
QjsKRv92plzjokNxxwTk+xXoUeKCZ1PpWgKw7OgZFeyl4nA9vlBj66SHZt9UtXkJjb5ipMsFugC9
an3bIbnIaXLFH/DXKCRcQa/OVGf4IknSXvLOPHX7cKZFBpcBQphTipO94FMOYdRS8Np299F6UgrZ
9BPcEafLvA86wAC0y9Q+GW/xRTpokyvzCYMASdAXUQErQAiN/BUMrfTQl21sUutl/IQSioXa3dmL
AQBm3Kjmjrq0/90Pe85fI290vb/Azu1aTzURurSvZINt+275208//bS1cLptdzFEVESje7uY1pgW
toWgyAm/xq+qIbt2oOopDH6oqzvhlmiSfKzKMBEmLtdC71n4LpJWguvqFieB3d6pIIP4S8KNbuy/
ajpxficuIRE54vsFtkbHvlVooBg6NxmPpguoNanvAMr0eESKmL/+Eq1UjZEhrRkyDAYPHzj31eJW
CH/II/R6gJOAPMo/Nb97DIW++MyoSbV58HYSVENZloAqVkA/uJQotdYf6ANuIRIWUmjvrFxv9UDS
nYk09xOnxEOVYGyV4CS9IPNBXX8QsUl9ef84b1Jew3g5kwKCpVfbiapUfcw2Gh9d73mRt1pzWj7O
ZNNPdkieXMM3bhYjKWWo3+IOCEDPKXQSsF0+aawWS8DnOBKhu6PtMUrhOpPw9LbQ0AlYVMOMNlJR
jE4SmPnYFQ5my8c84oMoXFS39Zxt1SiRQq5mxoWeHDhW8phv7F/W3ii+t8QmyNN6MbdsjOnNnbKt
m57X68ekGq2+m9NbE+D4U9csNkO2heplJTJz6zEtqY7xnvvC5r97Mk04n40m3UGDkz+NRZIgdJry
HuN9b0oGgo9s0Lhau5CTlxXHhjJYvGL9pZZB0rZvtss8TYxSZwpkxzP3/HNCH9K5RlaQyQckyC62
tYIfBzaPLMh0RE8nirJJ+zz64vIUEjVMGEJL5k0PuDl9sFBPKdovI63VD8nwUEHr8lkB96Kk6sRa
jj9bN8U0ZhM2JkvmC/aycuDF268py6c82opa2azmbf0osMuLJL8FroZerw/7e2VSlwF1mSF/PIt4
1OfZ01JaTlsF3NRPIbM+4zVhlP4veeFnpcALwFro9GnBeHscVZEDcb9o1G52P7tMY8AdtV0rHdjs
Rtij0p7hfCEDcGZQV8ZqZP9B7CWFy5g0BsbBPJRsDyIw23Ssynp7ROF21keJW17a1yU6XYTZZogb
FQfIsGWXl73+SdQnZjKBL/EnTtk/rwxC1lZ3fTXekudg/GI08i+VY6Y/a5CtgM9UHOvSUpPL1+ZX
rhOt1LblMhaG8SHPYgv3VokCJwINTCLr5UmZbanfYPa2XtpAxEkRedsvxY9cPHLNuq/6FwDx8AS9
fLEdeS5maTw943Oo4wwKVCFFrnW1MrJBNXXqk9ZdqSKcFnWdZ/BeWLCa83bbTYKUpUO90UJbzS+z
YjiJw7lkvOo8Jasm827CHBEKBoBFM8vvV80ZsE2zevke8rXTUdzfQVM0afAem6+PH1LDtDz9HUJB
5ljEybWFLQB1KXy21oDjfI4NmoFUutseT4t+v3uhXbBcQ8lwRAnhyj7YfDxOjSPojONKoRQmGiHk
JRmjtNL+AAJTmYAI91E0iKBUDtho6wc2PonRShFOv6vQceXlZqKyh7avRg+ZUAuo5WZ/hX8QnSeM
LdWztv5lqeblzflUwSTCsorFus0mH/kUW9dBJvJQ3p2litUGwatGIAzGSQsEhCRB3acM9Qsfu+N8
25AX3aKRYo8kU+D3eDfJY3OTTCvDrUVv7b7rnCKUsH/QW52oqzSJX8Q+cGyZSBuU134NmZSciIwp
TZ11aSd7Wg0cCrQbD10V3z15SXdWpFGBwRvlJhqx7xStOnvHbNForKycuiaXQx5s5OUXrbsvb9Zn
WYY/9SQQbi6xSlancISDfUUH0N6q6GPCpUw3dtNQZxAIqkqmL+OegnK2hqWsMcnsz3ByAJ+Ls3aZ
Szmh2Wm1N5yBobr/ICX2MB0v1SM5ME94/6lYFzOkdtsBZP3cvXBj+I1VvImvUJuF0YW1K4DTbuuR
ZZ6GpZ+xix+BlzMX3LruSimyCHoTpMW0Wf18Ygz4Wl7uC2pgwWUM5AAS0YdNvATL3bjAM6XwCHnK
6EN8jUQbdbLhcjiqQJW7lEWPJaZWBug1gsoff8icSe6n7JaHE2KWG9ED7se5l0UKvWApBRxPVCAE
eYBtLNnGMAFLeyUqCQqFs0lac/QQYgSI5caMSegOAJaNJUIj/b1O3WNy/oVTDcU+quSeqmvRUbO0
ioV2I3GSy7eAZxqj5Xtse0nzs7h/9MVT6p+uapi9pUHbqoGO1nNuDpz/nqaLYP8Q3fSNqCBvVGSx
SudNMSAdWEVycslpbsKDMrp+vMFJLQX4xEr5j1j7/R+2n7ZQ9tGC/BHVlsIw5KMHkWzHEZRHaDkO
tU3elDyV6VFdJlhvJoJ/4eP4QN9Vv65uL4Z4Vro+OBkJ7naaFm/BimFf9Jrp7MqRRbKhSow2lu5R
t54tzEoS04fhQnJogJyWnD/Dw6BrIuprmHmYH+CivK0Q0OpCMpVsclIrPjbTErdDH79AknFb7R42
TF69WLltWUunsRvPHwRQmssp8I4wi0fGuvdYVerMv3r0iwqvjfUZzsAxWqgF0GO33kgtbfLkf3a1
ku3FBxK2y8hV2fBN1mc8jMUbVZz66CaxRWucl3Dl+OXBf5LOPkpeVLFutrRzLVfVt71Z9vN7//hV
fJDwn9NMT7YIBELHXWIIf3GBpT6oua7WAzylBrUkAjy9W3FeHspMDL/LoEO6xQk1hLWcLXL349Fu
8UfX7ILSbz+xHtbxc4nPKGwd1prVvJQxPAoM2XPXaC4voraqLDSdjN1ENR67NAhNXaeSuqNSn/Uv
BxQRSv7zmiKnZDIslpJ7PR99DKroltEThAEBDb8sP38gfzGvy2/gqCjoAH1T050FM2CHLnJ7F3Ql
esWbsR74TCQ88GSkpFjVVVEFhkXsK4IX4ASBuISYEGL0oQJ7OAR1Qaauqh3OPUnMR5Rm85FYjT9i
fdO59RJG7QXf2BNeQfTiwfqwX7AVFJV4tuWGdGcIWc0Q9PjIMvx+lQ+XJGAZIt5yenUgbVN44XWY
tg+2FHBRNHd/X9kJu2en6Q//2ErsoNDelvYRNNru6tBKEGxYfQ61Tm2e2pBBDK/uMTPICeFbYtaE
xRFIaSPf4wIZl/Y43Bx5o6UMTrwim8vT5YYDYcGmhk10ky2JlAEIBr35+08WUSd6krr+ICx67pVQ
8d6ErMOxpi4e9rfKrwUWU5Zwq82gnc7Ff+DGf493H0H+VCKLSRR8SV7Vykpmx5quJSzEG+WXL6au
w/ICmGANT9ZRmeAPjTo6dmCxk2rq/VWpmzUMg/qWf5wwG2ebqbBIZW2KdvfgxZ0e+rdiFB31D1YJ
5gH5HQA2QCOe8oZ8pe+hD9E9t/JaqlErecZTUjjKGwVPu5eVmCFeHHR2J/YVXJMPrAPRjPBRqRA+
oUivA2iuyyz8/QooBWjHRbs6G7AKZhuDVlao6ElksHOYCNuBoS5G62BhWQ0yShEaD23NuFcbpzoQ
PS/871Cyi32CubRJEPzBMjskE6W6aYK0AiqID/RCD+3qE/Sjle2AgXsojEsoEq5hqobS++oLKKnj
uQIaNQWgbEtqLGXdVCrvP8D8S7Lndu5Qs2seZo+ucA8zkAtadkKmyxiBAcKunxyMs+7sHZuxCZg/
/6dIsnzC5w90oc+sNOQgFEtUXSJWtE8/p+rzYumfJq4n3Hz2GUuZzYYcWt2UKS3D519jORGjchGD
jUoWeG/AESh4WoAk4Pd3BkG78kZiPXskQNY2+6nkh80rRdGnLna0MAssm4DzM2yTGFUhtGElw4k+
aGrhyzYMYZm7y3+IAQyldRts6vpA2aDntMRTsUHTutWj24XsuTButuHIgzoRcr356hdRiRexnrZ1
DCSqV59bKNsedbgsecqaUFfiBqAUSZE58eoxxlb/qQ86IgxveGWc2ZJCkMxKrU6fulR+pXrDO4so
6xBbBT0eD4N8jl9pWy8TykYVJiF72CEgLysmo2QIkdJSYOeCA60AE7Xonk+zBzUPNI3ViNsjydYA
pG5OBed9EMADWYSOXUsNIJZ1MXZW7jbTd8xVAxE0ZQnsb6bQhTtv5k4lQ6JZpIbJ5CcaXQEtponj
J9f5Yu7KMqszWtMZvYWqQYS0BkWldLOqcfx5Kqm0ZMoa4umnPo574Y9Z0TNae5V/BNYjFdisFNDc
pyuE0tg8+S10wSXo7qctr9R6jHDkDK8j+1l6aWZKjRtuS5j6r+fFUqpLHlIgW/iazsJc4/nI/hBd
9sMOxj1LKTPNAjgAxVjvI/2izWoFd0l/TKxXhWT7FVeDTTf3LJsymj3q3m7ukowuy9eWRZP9PWUo
TXK0+UlK5JaBA7S6PIn6NhNjo0869uLx9uL+vFnVM5c1Ngfa8apvc0xaniRX+pIpcEThkdMWKwQD
uaqk8r5tzqOI1hLqtLCmCFoc5+tBbBeVUcPIaBYgSGK5uf7vZsnGUzvBe9exoSa3ZQhi7SFBTSOf
W/tgUqiz9kXyA9QL/SDwU/w0sN5avacTnafGUhdJmTRid6kA3caWPdw1kSk2el67do3lxuUZUqse
qBSSbXEgv1HE+dL9DTpgF3RE3jk7MqkbUipdk1xR3Mkt1oxqBrOY0Pb7TdV+Qs01BafE9JeWk0bL
e0ZnAja5KhfOf5H5+G8bxcmaPNB0H3cxHFXKSDcFm9T2qXv+FSCRR0Ib1ssaiMeKf46YduQ8MW9I
K1ZK9N2wXylriXPvyhHaE6CL2fN7UtOfvhHxsDlU3J1wFZPlE5oWarFTFSR357K/CDRaH+GLeoF1
tGgtDwF/cQVRfVXgjbvNAKR7sGlmp/S5nIDCVSzPoao0c04Yfd0XPWg3/EiM/824DTvShj1v3NMZ
PcwnlgQCF7Py3hNnF5K6Vs96URhsXVPIzhCBqRhKC+LyzXLFypYj+FC2xxrBuFPJdznJiV4saHJh
MUEbYvfHrXAR23JLGQJ3q9j7gTv6N/ZshOKCnxeHtkhnOw8Z0xMFQmT9u+SVBih5FUjXz8RdG/rp
vEtZHV6xqnDh8YLReqyLIrYHwYxMxWqdP9WYquFW6c9xGA9+Q8+eAw8U0kWykaSmQqipW/iu2Lb4
czQ6bU+sTrZTYI8hjI69CsRNBN3APkWypOQeUN/wjMoXDROwu2MSHBxODADVG8ep70yFGD9abopz
S+9yIK5Fle3ihRsrYzO4xVG9vFOlbSDlHeSR8Zi+94EQW0F2j0mLOnwdm9aI4uZhshFngzuNAuBU
M/GxEWp3U6IB0abLhj8A4MWAS2XzLm9P9gtkBY7uVDJ4eb9/3po8Tf58Z4fXhvPBdlKn+Pc3uhGg
wDAs0bP5eOiwTbmgl6Hef5ZC53+bFreyKybXyCKp4/hU7KigBVmy7hrZRMFS/27foWRQTpruS5pf
f6orvlYfzDyXpF1BiSEsCrGQWjauBh3HwHxC9ysE4TEZ+ahg0Z3RySZZtg6/MzplKztF9RJIM/hH
lUeO0Hg9c/RNc2dnH3ZwcAm85stvnoKH6lmR+jiotxkIbdWFazMxDqS3yzui7QNJxLczGVIOGCnk
bU5w7ov86qukOy4F0JuYv5Z/Lnx5UmCopxSGdjJDEDXaSxWJKDnIliwBgCuulGC7W0K1ieB1d/5k
ktG3KTgrDWkPlOsYFxEhq7L29rzx10BaXXdGP4kiP4PTzBfdDmB4hNM8J3/8LqnfA7LtFJLGq2RS
X1QESTMiy7GqtEh398SYUkYHKZzEaTerwf7AtF7wJreTaiOZBMWtPxhsCIsMtIGJi5bEObk0EMVv
7AmTu1zSePRKsLNfD6I6q/Z73OMqkI/DJ+vtNR92HpjTi8CFFm1DVNhqBdAF/vZWr8WgF4zVZqDS
Gi9V19E0ggQfsDwVVOGP0hp1YXs1hrWUZoJCJO9hj72HIGFbIkC0aDfjH3za+fZepdoGMcXCKlKF
WMwpWMzGVGn81dfrs+8vlbskluwHBhGYrIA9j7tzccStMnwfwUgoNocjgY1wbbEa8D2xudNg4Ln1
X4niIB7d86LcYKZLdQfvOXGEDFcSA6g9OHF3coIVr2fw7MK5c5Ernqj1caQycRppwL9lk8nZaA8n
Al+0B6wD9vqTQIFD8qEiUP3oApBA9tycRkG12iQu6w7eT1x16AvxraPT5O6aA8eY1i3hl6n2xFrz
bC+8wA/nPNC3e7j+K9jShAyYxRkp8u937E7ePIkn2bEeZ+KUFd0/hYxTZxgxLN+heumzLCPogGGx
Uesfch/GplF0yabw1Us2D0IZXt1oo2kGvp48BpEfqCnH9ASPxstw6OaK1dldYVsBe/Ab1ynynohg
Tu0HFY04mJbTX3JqVs24AXhXVXj6/8iatW9Y0NIjEMpTevAqEsTqrH7UFHZ8Num5Aa87TzHsW+/S
ifuQDGaPdoW2J6M5JhS4orKwXBieekyb3rdqsXrPtqNJdkaKwIrszm5rQBKKnI380kG1C6MRNuvR
5BxLeP4NVE96tB46J4ogQh2WDSAJPwnhZnbZ7kqHyAXzw8CS5p31CQ3jLd3y0k+06qGaBBW3eIMq
HgzgDDtmxY6T3Z3mYUnqhPQGS0PKmu639nXejK/xn6X4CZ21BJ7FeekpMkhkfwGiblAZnC6ndDk+
b+9KKNg5HaKc9CG4jIo3p9+Cl3+eFSnjClhfnUxJqoe7OEl7f6VAD8GPmai/l5eNx0AV+lV3PmXo
bB+vP507pu7AdyI3Xag80JqWaNi1ZGrVdj2srZO6kmrv8XXMIbAJLChGr4/Wv1bHG96TejCQyD0/
YZKhat6HKM8P0RqoX9nqIhGvdWbW0HXktVzpfUM+SOp63pS/fEMUSm7DjwVgHLO5sHG6Jt8wufBz
qZmE3520U2HDaJwkgi8wT7/M91Pcdb+2jzhlOnJ1sI15+jVLDPIxwZXvayiCyMXkgR7LAfDx5FyJ
aj/yRWGyoUzvZk/b3hR1POlQTic6xT+EWQRknvOpuq3ynh+P+8shHGMr74turTMRyOfFR0rcJyxi
EJvHZqkrm3HDe+6h9XvVJQuHxQwpIOmrzBZdMb2eypUGWCid1ii0lrGU+w3x8DrWRjQh3bTQL7pK
c12yp79an2TmxB/u044V+ggtcehJXw72h31HHczlquc0jyynBE0PG6gLLnr6+g+OGox1R5Piu+nj
bFNcnvV5C+nH5mLO8FhCj0PEooVerlEJ21KykXpL8//7dW1u0f4b9qz2opIKKyC9iPI5up4RoXya
BBUxVSOIFHAj4NB6o/UCsTMZmzTFnvPrAZ5ckiKMpSekkpaSO3xjVDGbOmv9+2RCnUaGscj/M4zB
NY+QulUJ5YRZaGkokTypHF5Xfn8XIQgpEKShMii+Q3PONWxQL8/UUjywZM3yvkgFVf+dE6Qv6fgt
IoUaBLqGfSlQWzy+5b7E8U1z3nX9UjpUnoavdNuL14wlQXvF6znq+HriFs74a1g06kSQXGOESFT4
G4VTmv+/wnPrn063Ih6mEnfgiQWsulzyvGUyXqYKgs2vn3WeJS9uidMXX+STe8Of40Dv1E0GvtaA
q0B3q9dHJidfiqTa11RJcJtXsrSH0C+o7JpP+TQ8PbJilGPQqXLokTM84y/CbMsSFI+CIj1eD5kR
lR4Efted6hgML28bCtQPqZsIdIkNXcdnB6kE1kYbFWj6lM382YvL35dLPu0IAZRh+kXVNFMNsIN7
pvFjU/T/PA/wjABiPb9XxkGBW3ZXDJr1E/A5W4y0NPc26z2TQqlHI3oZ3NXBu0C+Yp676pAC2ODy
yZh9wpLf7/6HdQKyQ5VYwWe0QKmrmc5oW7mGLGZ8Fo4X1YbM/HGT9vrP1rwoKr0JwhXz9ddvvvZM
YMzoyXvMMDqXymjOZLOZU/McWUGjSx9GD3O54UbjkoSd4Rdl1gh4eHu6x5QgC+oJpX8D8Y7i4vYd
4ZA+i/ldrhJsYUCVYCIqJo1D6X95igqGwbD6jeCiCwxTL507IMBGiTwsTbJ0NEdYDAYoP4GtAae+
TV0Ow89xnPkDgkiQ6eKyPvNxvqWjYBLOwKnx05HDIUrFPW5JkTemuHa1Eb3Nrj/pfnDpY2BOx+vE
z2tlmP5MAXNGEoOu9/PECLeitjalg1HLqqo2qQsh26TjK+ItqfQUDXWvgqR+gWpSvA+1moDQmyrQ
NaphB6Jnk+Kcw0upbRkTRRd2Q09Afz1PvjSY4IZ2/uXTAMiuyQnP1VCE3EhubTGJoy+QkL0OMdWw
5Yajj2FZ6lG/L1yGE0XXcZFPoOCDPbv3FdsJoKbzSIM/yuDu37TCzAryx8z1UJ8TK2CYtTzxQ/0k
VR1lfDO9wlEwMnSmCl0NrQbh4tuX2Rodt9e4d3kcG202xc88el1I4rpSLH75Fd8O9aSqqnqpFWaE
xgamdATopik9wOYNqLheyDM5MDoPG1Z2vUj+WB6TkjurPVW8TMieKy9PDvvPIcPVu0HuuRz5IA6s
LxsHXEhMLnbhBP+2IP91R0QmslpjpNnTOCG9jKgFO43PxxaI/+WwaZiAqwpNNS+jxDqZc2/elIl0
dAM3HLOqlsGpJyIGbs4oJ2vZjDFzTkeuuwp/jZQpcPJla4ycJ/t2yKSRyE07SbBXqbGdmw4D76G8
bk7Klsr4tHQ6sI1BKXPynlTtIxIVzpC+WLLX1IyYNNd4r4AAcoElz9EOzvxWa3yncWD+UMX5a5qg
qtk247oLcBcJqqyRtbwbJ0gH0nkU01aAT/NoOVkBXOT28RU5mshH/l3n46bk2aJbJJXzqkYrBNhG
M8yd6l4il42R9+nMS574Oor/wcSog6j13q+HrDNvYEizVVvLimNVCmT4CMzwOsBuuk2PjR77gURl
jcKmozub7z5v/NqXMaPnYELHP5Dn+uCNwU/RiFVlIAE8RNHFtdXfDD5aGpFaNe8e1Vf37kgDdIo9
IjJPW1mJcRUTSgnbRSFOC0pQxLg+s+zHp6yGkdTPCRI3bfB5BHO1xbsEyt6+RdqvJznCn26fPgmI
vlviWBmluFqtHydczVvjLdbzF0ab9o2X5BjlCy+ehUhPS72rBNf78HY5riD8cTkJ3GaOvDBngUiJ
wjor/Pau+IqSXGg2hpa8p9H1Wggg4XalIU0mTsGOZX9kmDsWlcHqeSvtiMuazPdwQ+C/O9hOkuD9
GIIJiEo9o1IhDwg2E0z3cN1oXvp8Zfs/aTqcI5wLo9SHV+Rv3XMkE2jmihPnaHaQfwYrgWBu7Jo0
MKfB5vOTLrl9tJH30AMHKBlZMXAARoJc9MstIbsods44/DRo12Z2+KGYDKQxSJpWvkvSLgQXdrBt
BSrB9pt1+POdTrXcKIKkLSKq+xSHjdAA2wd6GAZhc0hV4XzvneJ9Y+4OVxfUjV0CLrmn1r7kHZN9
Wko5hoGneyRT5WaHVzqJReRadYEx9B4wPrqXySRMcXLzO9+6CFUVam46wppwLaESGoOJPsnp7Sib
PDhoaUAEcZaioqqxBv5ZPgS6cOghqZXIzzU6o+smczM4LzjS5ZzMk+42mwC5NjeV5EBr79uYZ7t/
LJzubMN7xvUg9WCUm5Fd6rPlTQJs99UHh4vmIKGf0n68ozJ+BeeAZkqXvHYMqX1xcg7xz2+l1fJ0
AjK0T8X7opV5iIDB9Zioveq5/RY1Pv2PCV2uY8mUQ9+O7wRDV66+8oJfaFL4exDi3ig8fz2sKNXW
O0xKesXRi13L7HsDI8htggSg+5OzK5CFeogfGJT5kt1AfajNyJNBrYLCefgxeznF2Fm1y45glivZ
HvtDJrqw7R4JBVrKqpPJNguQwerAOS8oa3904IblZGS5nbLI+W2NvMMXAV7/PwkZ/aXeLN9bHL41
+UErNZLeOQ6E60T4IIf2WvXhIsyHYT2iddo3u0f6XgTXzBuojLbjASM1kRDaa/EEL++1+PKYzX6P
s75TP3poPxVJ9SU2gXMAnkmCwSi8J73RRdettQyOqesLteP9L70/+VEfL2IsH/Gdk6DBepGhnjTr
B6d29NLLTQeC78xGNdVNaOb4S9JOUu6vmPo3BfU4mxRA8elI2QPRC0KpsgAV6qijUa91Xcz8eET5
qwSKLCPcF7wEmgx/TR3ZLLYhHDVG+zPDqK93aWn5nSzxTzcF/zSDc5ysQQtqGLzkHvrCKHPcCrCS
W//ls43hB/ywB6A3TKFkTEMQsOaovAPoJq7c6y1feDcWzOusUIzgQuUK/k56xglpb5q7qlBAsLiF
9aj/GMNXjmox8N5rXAKd38utUdkghMSOybCCmUKqttcPz+cSCwJnF4Z5L4PszpBk5QnY1HoydJZ5
cc8Uf3boa6LeJiv3KQRGGk28rFoUm+xwKzjaJekfCHaLexusLvX6SxCS9aXpROZPWVnLsu315BIo
Gfz5hFM1wZ/QqY3R7mgH8Sfp6V2i8xuIU1vUvqjqCB6x6aZgDPXsjvqHxBNfNZz2RkdZ6PqbMWwf
AoPM4hs7Jr6pWWYwh+lAdj7lKF5XRQBmuLSyXCGO9gyKYaeigagFv+mIV6yJrsWdcEa/0+YoEVGX
lah5i0Jx/X7x22f9WBQ0s7mM+CF3c/K4ZdB6Bhlsz3c5njOhy2KNifilf68EOfs1cK/t50ZAzo57
1c+bGz5Dc8MCZXEigMlQRuTBfaBmnHh7puMI5d+XXs5zRbr4fPs/lnVxd3qxoexClSNWy7I8XqAt
wrVqvLBIbSD6oB+Z/RpRQNyxY3X49mlxitKXAbeKujHK9tUse+HJsuZIIryb5wWOQZIZHfppVSre
lAiS4jujMJkZYSMH/VSsVmt8+r3LJHmUY2Vn69QJdTgg0q4hln3v48GYdsi//vRipOMFMX7oNlEE
i8WYnu33NlRcm5/vA4k0FXChlxQVRSSVrzo3kWz1bm1AdGr8b6reQrQWtPNMgt1JWMYR158fqLCO
Gr0pMsW0GSWDJpDc7Oc6x9in3Hf2I6y0mTDBmgDTbUUoprXTg1ZTkhDEAL10zI80h6JmryiOXCg7
oW48Fs83zLo42sjeU8TRIPhAkXlXiAqTZGI2KF8PmZynn6fzDgahE3A1Rj4uI5e3aJL1f4QjtuST
18kpjxfReN1hJgS7wrQ+9VVyrFLFhN8lUgL05sEeDMDrbFm9zo0moUotfB1KpUF9LY0F915ICN+f
zpQxRQOsyAKlgSWb9G1p2ZISmpH+0DrTz5b1qeN2PVGcCv1BfdyN+Xpw60IQvbgEYYhw+EPA2odp
Tu/CVKJkdYwq6bd95MPiVxx2c4Ql1h+Gv/v6Q+EoQ311XoV0ppM5OZH+uWdY8jPK8nSD3Yb6ZrMT
6tuXRbtdzRyYBQQtPn0jo9kk9Z99fbo8ZbTs+uvEcJApMHn4BD5mGvZYQ5AAbz3U35mZwC0hm/sr
UApmYaKNXaOKrMBRl3vziZAPd5mIgJtsED7vTQIZY0mxDmKMN1R4k29mBwa1nlxYZlogMAPFBoqi
UYie5jGgYH96SNAoLDp0BDbZoV0kkKQiFpSlxfH87eYD1qIpvViX7KAyuQ3UB7QmKwyBf+PKTFL5
NkcU98MGNSq41M6EKZDM6zzpurUXQNfp7MIwqr46FvPTRpsknb+wTtxCSXp9JUAglTBBQQO6lz8+
nEUqCe46ZuUpXyh3Rivcvx3wOwXTOCLHiHE343O7+1u97lrVEuvQTIv7bMvFjwKWDGH872JXZogx
pN8sD/6XJm87tIvTZG7kF+vW17sALIqdWVOjCO1Dl7uOL85WW6bLShTkVpE11LMBbBb5axc1lmDV
BwEKgEv5sJdZWtco3czljEP9gW3Fu0z3uqYuFOgUh3DGyrcXcnKvUpV11zTSLMKDZLRxi3FV70LI
kTEYjzAJ44VbmhdWXZFSvZV3hfh18tKOWNpmkC4I3nCl/0zs6QxrSw8rf59wqrmMSf5EUfpwUJ+Z
jq+Wfx5MVLtBNdv/9vaGYFXB1ViYfEWC58WKEc2SqPqKmOzr41Loef01T7aSUhPpLbdHDk7dICN0
UWjcsRg2XiONS6OJivstFGL6bccPnqIvA//gDlikEUKZ356fJTWsoeMsEhwxI/i8WJ0zLVNjKB0m
rXlJphymIdAHZc8t+WxkP8ui06qDJWE9sbgtHDfTc2StA7E6MgLFCrYZ59Dfu1NHIdXveizdDw8O
+O3uzRvaJ/Nke7OYuCvcFDwg96zR+24ucw8ipcRUjCoH89JZuo/drAZ6Z2xx7UBi/+TciGARZ7Ir
iQDza9Uu4AYfhYNo2YCLlRPYEhpAaofZHZsR/J/HP4+bNvcCgoLlbMuD1m8ELIPbB8HE46ACqpzx
E6zM2NUI415WsyM5pho7SbiUqSRsnVEBoQmmUJGUcDTYV2qJIMoEKzs0WAjgfE7ABum5Sp5G1y7F
q2lBUk8a1AcUluaVvWdqmffFbUhj1dk5HwEWqBaMZrjlaqMKsPNktOuy2aEiOSApxRoG9afGMoBc
ITyxi7bW4b1G7hWYZipg11CSh5+Xa21BKAr4yOZ6udc2628O/PkQB+B8OP1Ct/gYbGSYjmZ8S/+Z
CVkyJ+4SeYhZV3NUZM0LTyHfS+DNKJr/r6P+a3avJs0Y0IBXoCr8my6fy51a4dSDgvdIkd/X/ZZt
13m4/IOcMzxo1e3f/Ipd8xnMiWNwkZFhMyheAiSy+0fCNqk2XDh4GymTYvn3GTjBecEroqWOeYR+
bkjt2KPjUH1qkZYBLFwTEigGDAeWznAFmSz3eAxJxcSP2s02c+iRPLPX8YZKJkFI82kU4vSVFMbx
mMJrhYHY+Pd5oV9BgWF+/GPPrvwcIH6ED7ZDl53pFsbk8p6o8uA3z2pY/xGwjdnohga58wfN3TbD
EyCXc4kGlbMFlqU/yBZYz/f60UawjrTgOLTLcLvn/0wQ7Vph7+AfrwaUZfSbvwT33lUNQpXGWbet
Ua9/+Y1WR3QXa3X+TxbG23TOhCoCrtVDv+CVmgIPBrF8576bRG0I5ewYAGkqyw0TcstSJT23YDXY
+lknZC1bw5uBQ7v+RSOV99CK1sOHNe8MfAy645YZoj/E9a6Y0zQfc5AyGswZtl0peYMavi8/90ji
hwHzF5HDyEP0iTeqH4KHMnhoHElWWSWaboF9Ke3o4WupOT2eNXwdGMNo4iZB8/cszd36kNP7eEvm
DS931a8cb6jup5/hLw3aaksJAtTDYITmtRQxrUxeKuAaO4m5CYELvR1JwgXelmGrz0aMKdWEUtfV
G0XPRSrEm2ZYkeo+QQiLub6ePQ1keN5cgwFHogQ/7ltV2hDcWzcq802xqiR610EqAhK6Zw/XNI+w
8iac8rxQpaNp7T90AxBEgTf4FF8iCuRcHxtD1+Z0u7QTHUb8gN3UOeoEQy3mfoT37o2DDEGp1QGW
uwh5KHhhJ5j30/4IvkPB8lcdc8SG5o3L0sQWssNpshNOVpXyZh7/Va5dg9kQ6eaCRiDkvpFvRUik
gD4TcAOOGtQ5W1+GJcNwgLcPX9zq7txLQoM+pLWs6fm2wUigD5KduVOObHvi0XeEeQ7xBCuEG5d1
ZaHgwShO2Yef84fYq2+tBWleJu4h1NPKm6q3NOXK3UsYtIGei3N++YBjiLPhSqQL9RIvcs67ep3I
jMO3cVqexogZ+Tgddp6y+8aK3twDwlMPkrcJCJysDvrdHgVZo24Nw9w/bWphFroJOCLKoWT9vLcC
ktEJ3zYs6qp0p+VdDfkPp6U+KiIUHU0zT7gybNh/pvxh9grtMN+kY49OJbAiyaGU8B1C6cxP7tYZ
xT2tyahc19NpurGA0K/Cxzvbf+8fXFbXxSE885cq5tMHRpoBUz+BxaH9F8mSc6eEXyVnDsz9vDmU
+oU+fYcDOvTWG/3fBUANZ2UOCJfeTydRUwNLFveBS53j5vM/kMKr1PKZDynNhMBECeVaIWm0WF98
HwgcqssIZD7dRd7i1o1vj9HEpHIWr1XpSPOmGp1RyXGJlz9P1V+TZgl5l+kbtCLBeQ1ZBSBxLkZt
B+Lnbyy91jRdKEjpAwl2y8UgsaxaJth0rW4DH28mM+hMFKIwmGxBytj8I3iKN5grVc7DDqE8gmqg
fKTbhHBLKIrDahNQYX9EsecGzMddhVB37GjMgtxXUtXL6bN55/L0SGl2uaJl5FYP+YoO+6yXGlho
Llt/LeK0n1KweieNE+zwwhjIhPW7E2VUsO7PPOEGCAdx/L0aOuAvLszq7gGEVym4MjkTeMrnUBPA
59pMxdcYJe0i55I50PJsCcITHZq7LpPpb5c51ob6nYFfg8u5IMKDUKksilHtLGiO5qqYPTYoK7iA
1zN8J7HN22c0VFkeUQArEHN/M17uepLbUySX6Z7WoVo0KVcqBGzqgp90Fm8L3TD5Usl+sacp7x6D
UT7nEiDzIjXyHd+SMtAsqaXhQlPzE5KdrsnnHRDB5Al1sYfjShK44mUs/poOKet+voq8hOncJnKr
WpRYF4jdEuSFrx88kyqOvGkhOr8mcY2HOlQOmXio5JsiuZ+uN5wysrBnQqREA1S4R8r+7FA/7XG3
xmVutBjP6fNOcIq92sIEfsbZTuaSoGBswvrU6Syx5pK1XPLCv8ZY/AYQYG23nchcGFpR+NnnulL3
8WjD4j4g2hR3zN+Cs5EdXcx52LFozIFOrMRU6v2oNX7JSSyLSvqzFmkbBFi5No+zgs5Tg5JC+HoQ
rynEM0DPw97qSQt8KyUzQiU3RLoRxr9u1+L9y/M2n9uAD8EzpU146Ck9FSXUQknkgDgsqXWVTpAD
ZdnDlOaTUiVWHsibp5rpBNsz1CsaXXYuuzWc7nsDxOWakwmSSbeYjgGf9GKasFQEwQ6V5fQ/N4BL
7OfaPJDNVyQIVMn24IA1VBJ4l9yY1cW2aeudvIGZ5cmmPkmmUt4T0GUzHXJvv/jznucMQPpPMbOp
EgxJDt/50Cx6YySC/cpvlm/0rZLBPt/f2P7K3S7DyTZ8GJUkTVeh0M/gm2DLuk9npUoDoExYmNIJ
NXxmuI1voy68CE0yD36OuGI/wRGqOA5GcunmWs1W50NkXpsd/wAMZirQq5qz8hKbJW/eOwCgLrgM
tnMGXAO+XelG6lKwXuRmXgVEsLOn0+6dAKUgB54aTOm0WiIvjPlqVtot/ZsqpTjyy4HtiaQOpnvT
2OV3HNkSHdsA74zvcEXhK1A4O7rnP9RSdnIAWHhGVe+ekKgFlSDdAq2OvT5DdsQoatd7XaaOr0PM
wbEciHLpVR2zbmKWhdAwhsyRcXkWuIeOOudZypwKQJVPLJxa5LWK5/sCNtph9FGqJHMVK6UuJWzT
BOevUoqyS/Y6QmB6TLm2TaU37ri7J00knft23XCgYaP6Ej04zcClWQvXFkJOYva6c7TzSkwi87Ct
+e3omETXm0bIAld61gH5GazMnVJA3WR0UDLfCogbgFTNxlXQLFpGE3bpCRe4nF4mgaPLECeVdpAG
pReyIPFDjBspDDysUSj9WQIYmMZOFDY3y388uUmoWSML9uyidxHcsKTHs6SC+rZVCwKwPxacdLSX
2xjzhmf8V93Z8SzxsqHQwAzPoo77UDhrB3IBVkPk/lhIEEFGFvMKmgl/vpIPoKzEve/JWrlSAQh3
8Xt4IAyA1hoFx8LJ+89TZjudwpm8TNqhKJSP7VXZ0xSNjHSLOnu0/8Q6vfqC4vpxDaEeIj4sd3Cp
9TSTCm/SCcx8JLeFnzFTvFBwyo/XAwHGfAvQjgmvnJ8mL4k6h5BqlYy+foX3pVjBZSvy1s+sVSm8
Ni5Q0uMlS4Dop/wgqVpqKa+0Qk0ia3j8VuRYBIh1xGYi4/RMc2UDEJPs1o8yu/i5+JQ3nsCLQKzW
L8a6NiIIia2rJ1AwVQsoDucV7XuOCNPyv3Py/34bsSB/65D2LR2oEbV0KNPgAS5YwvZie0J2BWYt
ItP3dMRx8b7a2mzdXs36FMVi7dWwmXHCunqpDW6fHh7zJeJmxcXCNuw0LY65m2gdl0fctA6W1KE0
axDYNssP/QyAU1GDiE3bvCGoEixEjJcFnNbaxW2XA/Go/K4RSpi9koKWMRLpx3gI7c57tqG74U/3
p1rztPqcu/1AjV5tSK0+qmGlEInqT7BO9t+SsNEyySN1m9ixsFr1R1qhLDkLLPzkhjWcojQ8uLxh
GIfBRuk5DlU0S+TkVy1Lwucw2TtQqRbA6PCpqlIYGmMrI7PfAg5jVTZctdlyVqJMQvqT1ickRqdW
ImtMOtoBfKWVrAA4k6/WHDBUfMUUe5wRmsD4nTPB7ucM9YRfOc8Fuju4O2WEu48myxPxsJYKIiTh
UV0SHzt9aJPiqK9v207v3BI2NbYwhqryCU9xyUHsDNrmBz6Z5BurijJmnG1jOZZgMAKlJedbyfwX
TGxje4jmUBIFuXiZNzcPcTT3xakGHY84CvmqPRogrCZv0Z2KytNLEjTQHzc2BCuwu0Z5EK1Pd/nt
MWH9Rwx3Zqsb68NHUcW7qrCGL/MdCB7zNmq+gWEK1EJHummu22Jthc9+Qm4tejtZiT4EQPhhunJi
mWtcGvNAffO4ptwcIbKwbCABTK44iI+VLAkVYnU7wmqh+osOuYcVrQPggVGp4vEKtXcunhY2VXp0
pGgCoDaANLR5lowiH3rwVA0YQqM5AJtkj24kzLShcFepxu4XaTQ1TIqjrBjtuWsqkM4z1uXcosGR
4C/BieFN99EziOkoLmA60EBOCtqZbR9OJMm2SqTwpM5BjLemRjUuWrWMNgZcgH7xNlXDbhpAioq/
kwnnY17OX5JScD2SYseqierMHVSnkHr0MwOTKY+b3uveMMsZB1ensrnwRFC8ncPn/qNSmFPVNzy7
ULTvXWdyEx25shnfkhN69OC0qHHG+Le9ykJ/9sGk4kIutaX1H3ke8sOayyRnmbaGMMd5SkCvCsUp
id5IsPCJM1NwE4e6BhkPxOSymo4HnUxLxWAv0V1qbdNCvZZ9IBaeIiGBJVbaPaTAA3XdiuvD48vb
T+C8PzUaryixGQFdND06B+8fHIvUFSsIobYMfkfzxZ/kj4X8mwTTRzJg2IhmD9XFYTWLut8oPl5N
fuJs0yMTjmZIDKe7ZV+leSx0mLTXPVvzZr8z6YaSIv9rPfwW7rTVwmXSRzUCDOygoZ8JtO437ojA
Qqs7TlKDCZ1EgYSBYqv/W0ZOVGabo3fO+F/Rq4Yn1ZX0b3cZXvRvQDiFISLTFwyNMjM+ABUXgu3E
fSLl5lW/6AjPvY6bU0/GpVKnWQV+imsXtWLvPVbzrOQsu38fgFhGgBmgAFuy7Rq28lFxDy/uSb93
inKASHrW54znfVBO/SfdnEt5T4/m8rWWb0PuAc2eRh+GL0LmqiVSWy0LLB46+hC1FBOZ1txKXN1p
jZH2/Mhx0VK5Hu3BKPjuG6+vKIJCw8Qm5EAx68RJsUd1EGr1Xzcjn/UDpiflQqBrtER5aWiLY2lU
f6u2vDwuKQ6RgVT53IbUwCgNs4asWx1inBoozzlYga2/AOw0AdHSMnOUyMEyYSw7ecNCEYgJTXsq
HcDMM2HJy2/pMtQ2C8H10EUIP5cXNTaZkp4jJSenZlITDl2T3jWURKTzYSY5zYkYsofVo1sKIiJh
SxCkPSxgSoia0PiQO/b9NszEP7msCDHTN+9C/Xr0CHNvO3tReO/SL6tokyftc7IS8aXoYiqXQ76t
eYLaUPKZxkCAfvkKlduy0+MH3/rOnlAqFbj3QzaRyw0mQJbBl0H6afbyUiJQGYbDb8B0Dwl7B+13
1vVg+Os80fxTERct5maLmYNqs4K9eT3OzYQ1jeIM349OxWAUWWBYg4Ua1smFM84ybrUNNeeiAkcs
Y7u9qk0FD1v4poYrc47qf+cqKWo/qvi+fi8PPpM1x7G2Zi/v+8+QcLmR4dfSp5iqTSuWbPrhNG1N
G9NZcWyJUNAeun1tYXoRp3Oz/rXKvj2tkIars8Hxc581iEY/u0BbJtlOxyfW7WUunff+8LVBQAWu
oka/UMxvnAIGWKkwcCLJZDr+lxqFMMnFolz6T9HihdlNeOh01xp36/5zTi27YRqfDZHd7IkdA/V3
hCpyTsF6twjcFgrotI8xBCMDIJHDx5ia2sUaASrAEfaKHqpIj7zMXzlUShUPvWbm1f9Jd5UNdiN/
hgHF1iGtCt/fyotPZnWyobRarsag8RN5tprYtaUv1aAjxxL2WIOcrZvbkWXqx6AwGGB0qn8gvjHo
3RWr7jDElcLqUe3IbAlO/aGFwOzX25XI/lEbzJ+9FYbaRTzDC+dDn1TsHPG8QHqgvHIMLmb/6g8s
1TyVu2E3Q+xTFqn3zXxJ+KvBYMg+9OSlpuOF0td3vza6qVL9frOxgqw6tbq4DIW4h2FpHYLFxQa9
kJdbvsP8J/XJtvfSbOpzIRKTsuSoN9lvUxNpjoiEHCcO6zQDEELrNnnJ+oE3A0jd360cD4nG3jrf
6SfJok4uqp5Hd5zjASSjyn3dhZmfPSDYW+/+OLiKrSj+ftqtqgvMxLICbV1H891/oCUfMNxTtZnV
/QCFd3lcy+CEl2VlDhFT9Po+URwmw+7shMjqfxD0W/siyQ3wckXJl/QeB3snNg+ej4YL70oRQs2S
jQfxvkDIOlFUcCc7t4CRXvGOfMbU2Dwrj7hgAkCNi1XTPLVHv9HWgrRsKnpcuMPHVYf9WY3W+Cmu
yn4uM4xt52dFZBZPN9gB+Vji+jZ5382qF8lb5EOXgEwXfz4hPGD0vnRAz/daXy9GSC351IWBypms
ZMBwaX03Ph90GE5CC4ilsv/TXeYynG6ZCsIsOeXoqHgr8lYVcf+XTpu5HTQpP3aoYM2YDGjeUNl9
Jo7ETVTm/UjvDoplDPhf+Y++X49A1WGbOKNbvqUUHOsN+pV1OfTrccFD002FuIZ79WYqH4JWUUZT
EqO3OIR59WLe1fKhO+U9okwSccnooH5YQVyP/S0ocmj5OqDyHdfkumMC8jXXNx+m3T8dppVM3v91
/lHBRDNK954Q3wv3/Zu4IUXivNaQ6xpVXTX3YjYoGvkg58mK+C0XzO77QyUTWDygvh5oop++/HKe
ERYVgbV+fC6UHbuNKoqQiG2s0eq4E0f6ehmoIpcQc2CO34le+AHP6CrTP89eTsr+lLoCSBreIjbN
/SbSxTR+WUTbOaXtACD0eRNPE4enHsnXSCdxSWEWCaPuH0T3uG8CqrjdXwlHwBW1bqr4lbryhh1K
zcIP/l5LHqY2cY5cVPpCIUIsYmCRPZRPUUGc/JZWv4G431d/hiLQSeI7wY77AbXaBbA/uJICkENs
V9TD9kLiL1ChJDixx8FTKqOb2zJIbA+dwN5HjOCGQGy3oKbgvXZYwqF1UZ8OIPZSmG9XqCgEr5+b
L7QiLS7EulIQAx5PQKFZRdxRGF4N6pXFkBl1sqzikDPZCg5j45Z3QlUy1A8ABf/dFwQ6Ff4cmBjl
shZYuSb62whr5FIYOYRJI2x3hCQf3rYQmrm7ma8Q45MFbtYvzHmnT46mK3GIAiUNNbp+dZKeAUF6
EV8UkI34GZSir+S/KCZy5vQu8m142335YorW+DmO2PrZzNSkZWUBSAVZMfHTH4Qkrnj6rtnlDFPG
B2e/UmC2hFtNLc87rCdvXY3VlbIvCAf+sadOcv2CQ/En1j+1MVNMfG4Q8Miw8jCoc4ZY/Rd77WFW
C8Su+7QQegX9hfFUOTetMzs6jO0tKw55GXgPWskCdiNN6ASqq0+qMelR+CT1JGZpFa7Yt6PJpio6
fqFMO5My0ThHDHQsPPttFhmyhM2Miy/k8NLoFr45thggKDaozYcZlbdFH4Lgn5Yuue2Z5LS3u3wD
1wagZpgAnwaE6J3kjaFCDRyN560Lm1tixLrfxG5oxiyqpmtCronZf/OZLtor/eD5GrO9KqYyhWQ6
O+HZtYNXrNyMy4OoEOfaotDuh9FSAaTKWywAmpxPhlvw0CCuO/7UBYj3kAaP5VST0SXJUu5vstS9
e457m/QQNWk19Z7z0LZo7nAE0Kc89m1bKuWcXi/Szpom5xrO433iCJ9WGTCNCzwb+NrL5S43xtZ/
ByOBr2K1Sho2+uPVl3Mx1haXyRopKt/SqidXq92e5kTO+aa+y1Fk+6EuoAvtlw9OlUjIOUMFJDqL
vu2sHHyWE5NXRY0BUHhDV/RFqTZyQPFGzdzX+WlDsBsFoXWjM2EoFwJcZhndkc0iQdMV4t/VAqb9
k44DdA9ao3/UZFQh+zGUiWw7Z7aONzp1sIx/TWwBvMc3nFlk03DgNda0hpkIZXjuq4J3CEDnwbAt
xpdvBshnj9H02yM/RNMSQia+5DV5BmNjaDBd3sbhk5HaedbjKVtbzqIooulToSCayDOmGkULHy5w
SQRhyHt9Ck5miApz5zNkGSeEnHc4lEw9NLIn7Sm0brrw67UrHiFNhW5N3DMGYl0eOo2c0U+8UoOw
dQUjF/XzXTIdCo134XzdZ6PGiJ5lYM7PzIkxeIfdORDp1SoShMTIMaWCcVllmlVsoacY+QI8Svm+
r1sKbees1AMN3PA1g3l+/62wIq+284VAa6RZ8Tl4vrPVLagNtyJ/ieTd3HhuzB9nwCcM1Y7FiFEK
tm17bKyndAr+qYkKyRc2xar4cl7OMgWH9/RS2tGaMrUkwtIC3T5C4wEhdAaek6bf1BtsSNsyL/bS
f0JoNcowr0fehUc8p0RmS6GNWsVG1emCJRPKRG5OIMjF6tsPi2+zFSM6WT4DDL+9A8vZ0/itMRXA
gyuHzUguWtwHWN09ilNy1NwlvEkqanhwswoTFpBZPyQFcvHwMc+4cqtUbb5rDRU1j1EhUP+pBbeD
sUbWQgRLmbzfv14XiHGJRjYxliDx2/RswcY4JUtleMt9LrVpGBLsxp7xT8hYe1CByarXk0/C623w
edyZnF38uqm2U34NbhNuisc9cGbBYGM4l2Q2hTJ5IAD8VgV1xFP30TIPjbrjDyKsVZvp5WyxlqVE
BKhfKSosV2/bdfcBBvvAmQSobEE/Gw9E+uYjD3f7TqwXJ9RmUMYSeO3oIcK7tdgTEHjdSaCdBClW
dOnVWYso4MLBY84c9FyhsqDm2D8ia72nMWJXyP3Ld4X08lnBChUHDw3g2uae0z1j1IDQBvvmK9kK
+G7py5m0oGHXFjhVtO63KC0OQjEE7/LX/aaUEaFbhQwUsexk1x2JrTmd14M26pvKV6IPyomw6w2T
uDkAQfl5vVnyzJE8Tz3Cxhks4R5WbLTzE+7mdUmIGnNzJNw+Rb+i3KG0olv2Mkfg3n0u/3toxafG
py3VdvGaH3jQepx+WgehuwKb28ZwBhzrvrTbv7SthM09X4oTyIhSO6Ylx2q0JDEituUNblkszxrj
sKyhc9ZflJwdqnKTM1Y7viRrW+6q1NII+yji2QOZ+Pd0I5C2Ce7rgEh/zNwMikf3J6V4x6okpsOe
pyx4mglK+X69u5sOLMw+E9ECd0SGCN2JTzZkLqi9aewb9hmoghxoYkFA3NPclt9R3p4JUR8nKl+S
X3x31VFZanqjpOpX6ZN1hoZVj+EvRRLpdskutbos9T9QORJvomFYL/gsQxemQvChIjN8fCCkCugG
A1EyLxnbt6NWucMK8K7IX/LtyqMCmASYMkXYiI0d7KL5YpVEUWw0OOJoUlQL2Oxoijxi/+YLXgvU
VoVKBQnla9s1ezdF7Wj8vatqpSNyNRLOal8KRNrbhoJ4zquPRSdLidMGzD6Uis1Upj2M3Nfmspqi
uC3sA/nuEN/L0YQTotI1d0nk5LIGJbj33tWmvfQmxD230hlkr7FbW3EdIC8MTcvH/noM7/tkh75h
B1XYfbfRQGJuud6JeVobDUma4AYtgG1aZvBugrR+UAlSq7dsu16aeRMj30UT2yU93MpD1soFWlNY
/KMIkIYNbERvpAWwxOFyxMj30U7OY90gFe+5u+AKzhZFeX6et9Y+99oXK1LrvbEjCw2+p3bGz84d
jBWgKZlV0/F1fJV1c0nJ7Ef6vNch+DB5Dmdxpi7Dq7lzAS+uTsJ375EHKnbD8xpG2Qq9nCPAabZh
ZTzIAQoLB3KXKF4wiNUvvVwhzIA5TwZMz9IlWvAU7W2hezsiT8+xOg3QIfJsO7YsWqrEIa8jjg38
Dh4n0Yy4Ik3H4RN3740ynJy86UQGfr3hF/XZr3XkTnVMD/FO4/EvpS4BYzxuSo9xN3gF7F9Mj7xL
9sSuOfbISVMTZHJP6Q85qk6KimKZ+MqHQc6MX6QDPQM6tVv9zvZQNmKLS5mC3eainqi/QlwHEiBc
D8tHX29JwoPEhHwNhtAEYw22kDuyXhXvQBJQdbcBczuJVpvsy1jmdfP+fMU1BMvHoqQrQwdFjyHE
4/Ia/X6ezUWOyuqSHzaGFgxldibYPA==
`pragma protect end_protected
