// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Yn/xG312AZigPPsiW97fR+ESWphvlkcDyQxJZoCBdiyCmcHgWP3gyZvaDnWJgK/ihgntlkyCyXdR
zpAi5AGgMXw26J9XLte/xj5ba9XZvOWQcZwOKYkr9zD7n2Od6DK0J/tREpQyfCRjREBNRXkGScig
+EJliO1tBIyZZ7ETmIeMQe4KX8L0NsG2FDzwiBlLT1Y8ksEwiyIrn5JwgTo8iPPSnk1d4oXzX91D
/zZW7S2nf5DS0xKDbF6U5cg7ZCewdzXb3CdF6p/xmu2XEdjtY01XuzzZWzDtwvcqGPtCuzGMFBru
0VUnpXW7bEHw1QpRmhVaLGq/UN7Asb0j381Btw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
uLlqc3gdpwzdFsMV2a/0VjB7BOrgIuljLGoHfS11LqBR8chiz9kEV93Cmn6qsEXGNu4Jogi8lqM8
0fZIiUUpyc4+6vwgC+mSD6X57forIwyF3nI1FXLclks4hhTbPZgQvwiMwiVp5Qs0qQ6BDflB4pCQ
/z75p6Y8/4wqsR1gs8YPDveAf3smnbev4hKJ1vdswU9iJeiNK8StBc9EPziUgIpoF2/OTVf5+BZS
d1gMXJlEy4kk3Azn89YVpwjTHbqHhnb3DNJEf9THY6kPk+avpDk6p6zaOccC1riUY6HeuPWyBIn1
BiNo7PMfDH3/sBGbJoM/OIZh2WFhyuJ/9n8ma6qhwLPOyofj4GlSk/XtINlgLR2ppwyDCMXq39sZ
S2TvqGkaIibtT6tambbjeuz1ZrNdxiL6y05bBJGtVq5JnQRhqJFm3UPkvxLGiU6woeN2xVbPgoTw
yM9S8aPDoQ8WQibpb+vnTxOwT28ws8o18xv7Q92jMnbzhUi37/o0wNOIVvgF9tairT8P8zQQvx08
W+albvjv+oOepQQu4MH/qo1VOEU9S7TC80LGSjXg7LfuSUboWOBdpe7QDOrc9h+oY3VrmNgtnfVT
7VtmjRseNGRGAwy/vi6TYmh8ecX5MW/bqRDnHn1PPqdWGfDNsSdVeFM1KBP3iTgfUUgHZgYk11Jm
GSUDQO50nRUnijcpwJkt1S8+nG/6htTEanJWQ04awHRma0VCQkQblxoHDmxwbOiUPZ+69GcFpldj
+vo3HecNrCyUl/hE99f8SPzXFDUSmgnLBghRNEsljHEs7cvjCBlHh0v6P0rbdzRYE+KkX6XUWcDt
6LBqQJi9sYGqocBRfTZrh9g7q9KgMZoO3SugMDuiPaMO6TmAeiCJlNRAhWyOpMj3Lg2X+jAdrKYu
IW4uO2s1R5bRWQX+fOh6Kjsv2d/OFiOTON3hA19jOL5QyPuxP7zVmoiJFg9o1j7x6QVt7/H8UDKF
Fx26WvIxhVTnkzCUn54A20y25Rdw/texC0H5gPBvChzoHy7N+B93zn5BTwMwhSlYUZcoHcM/XzZm
fQWV+DtZRI4fKvfAx1nSQxJANlhU2hUSMhTXYKKZxSx+ywxdUcDZWx+lkLFMnrbIJ7lK5taJ0ZD6
MpvCIqIDCovGYlVLuut4AWSVUuQKcgdsaD67mRBn0bmXl7k72A+FuwuUS+RkwYIdbo0LqxXkMbMa
5ipp3HGVns4Jftz9Wvt0h+tc+9v0DrRtifFc+mBpHgv1CnuKxHlAeqQwxDAIa9hbn4mBT4kIn7ez
TGUGP1WkJLSR2eKNyv5vTQv9MD0Q5xaKYucz9lFzHqlIOiDq5Ohcx49RryfEO6G/+NkPh/lJpvui
tOOWJQmgitq+lL3YEgCbK2LpizmiVNuha3zRRUrN4aIxIE8HazDzMfyVpYXzOubp4w0kSoecK5KZ
w9q1S8xP5bwpWBhU5JwGagATak6xXRwxmdw3QTLvoHj9seUtEvYMARj0lVuckXtWeWOw7t46AsPz
zANHuBGi0UOm8hRHMd9yfY0cRmOeWoB+5j5jXwRGHiTkMsyZ/cJdEIE7iXmPDwaJIx/lEpfM4suZ
IRiTRipYD7sfUG+IjA+w4oxDH/4cOHMtFNKSC9Y8Px9IZff1ATSoOQB9uriL54dg4zgFjyC8qzHC
ezklse96hYxBQoE06CBXIQ6dY4BMStO5AzGrlUWtXRfJ7g0JxbaJnvNh/VrxmnMosNDjBy/YXxuY
llhiK0hHuAmSrl7CUHlJobzJRoSnlLNC+RCzov3Pb4H7/xjBVjzDON+EOBJE8OaecQ1zV9jS5m7+
pfFCXPKfLO+gpidQ/sZ9VGjEM8s6VWhw92Dh4/0/7efkeQS41Tl/pn5LJKsh1I7QeBwvv1xv/OeY
hViTvkaZpZdRxc/BH+xoBodMP84Mh3eQ2rT4/SY79z11MXgclBTpylCexmeL27lXWT0FRkmnhUQg
QbNMiuVCJIlclWNiPdAqNDAkym69SzzNMwO3gazQddExmiJ7T9E/zQDVQxSFH+5xmaoRh1fJeEeW
Y56be9jFjaEFcOFa0VjLkPWshm27RYVhB/lGeSDUWAgpibZtEz2OnYIeEPHgXfjG0D0yfO4jNV1E
32vWAKyw9Ot3fjj1fOh6ZmbMZM8IBdJpUZKKwMLWd7/fAD4NdftnADZ2DtOG3KUDmdAR95K04Tiz
LO2ZNb6aOaScr+5cRmVjHoCIKhbbYtfJMuiz6sf1ngWf5VzzYAM1DMvKoS1CAaQ23zrXysGfyFZd
9Ub1LXRZ/g7gCVh7bF9WliFJPWWL15Aa6uyzNo15KRGCstXVsZeyvPwbD2lFmKSp/sXFXGBk9lO5
NHuyHimJZi3jJr6h115ca+Pp5VZ46gA8Mq+w8QtQVrXtLX4HRRJh4TZRwT7chPfI4YlJDRW7i50X
YBwZfaHmlybVgzIKVV3wmR6CIqrWMvwRQXJieoKS+6DnSiH6El1ko8aiI4XOzGVMc6Rp3D+p5sms
W2r4Cabj5UhkjvCobtLaph3iguFq6wBXwDslwWqf/AU/X2TI80pWpiR+/lwNgqIGpKDBPdWGmeJQ
b0Yh/KKFKKzK9Qy8eSapFyoijwPK+xFwFawEfekNXky0tYh5KRacZbXpmy4QeOHaHDuYlL4rfogt
4C9vs4S6AEmI7ovuExtzatCs1Cbz96gm0Vf/3y/173j4Uu4k/FYYCHHmuEiWYXLnRUin5/0TV2f7
ZyNI6jE5v2fyivA8yOZcAXlmlDtvCMmXOoU6590zsf/K1fTyUucaT8ugEY+SWPlCPXjtYVyelFmH
YQskGe4C6vExij0P6y+MAO4oAjWgS5TWPkXzxz0BUoseoLq4w3OVCymcaP4XYFGRTafwlGsYJ/hH
xn27L5nSYamNA6MyeCxG29w4jpHgCGN+PbQPKwyeO5r8fyaG1b0oO1KEPVGHNmIP/p5jtjSpLNUS
DI0bVGqrgbYktbmSmRCEuIGfzF87l4c4/rXn0Hx5bcL81EdLrb8gCfqCG3q2c8t/suMr9yd01e9/
dfNSCcvhgb0M05gviVIJQS5qfhfuYoUN3FHgcl6XKo1IEP9emhyBIECGSm7oLtjQbxBTV3aMPiiI
o2F3r0KR2p3nH6gsuSlPnUaXBKxO+v+RTxohzvdaOLC2L0glJliCBDozoDYaCrnC84azuOD/zeF+
Z5zdDrxX0N2N38zFbgg+9W6EYY+ndIolcmborz00OcR/iCms6FU4MwOyS/mKpjB5XJsa8om8Wi3k
EhCd26ZqpbwI8YvNmYuHV6PkF1HxjvhIbISqJo8+lKyWGU7H1vajqmnQppL1VL9D4ZbUJwOPY/Sq
ndgREsNg9Cjvqw0QQB/jg6bm9iZl5uditGu2nZWArd/sfdLH4rjLnIkCvYM8PJ+UhRsEj8sRKi5z
nKM1k0+x481jzshiYe6iP6RUrGoCBlz10Md+nkNmvID0ZTnvbV6ZUYE65/amMYpr4THZzOet6V5g
MI+x/W0iwxDa1vZ7BWK9IWOo89l1HHr1OW4XDii2nfrGFq9WcwY/fHh6anAcl7fZiP85QQVpm+To
hyK5T+8Tcq/MG0r8wDWK6TQ+VylI7JrWbNiRW5Fr/druoCgb13ZO77yWiQeHORicRJyZkqIyLCgy
ACfIZzW7KpO+GaAx6NNOLNn3x0qONtbxLPu1vkumWVaK6zdLZeyhMOfEeWQzaub6fs1DvAPqsjDm
JQrC0STp+G3rq2szRoHCjiERsHo6wdynasohOcCYZpV2v6FpTs1NHesivfFy9jOboK9w24yS24tD
dd4aCNqO1ZJcfDL0N0+lFP1G1oX/VtC0FT8MZl0uaekpW0vMmWBhrapiVixC0xjrisCjFTlRFr2A
YVY95avXvTW1/IkRmZkzCUnTY93bZL2z/cPYZkMjyzAY9S+utz0ENReFUXIXGy7WznUyLrUSWMag
EDDkdSjdgPMG5NFPUPaNFkhngfcaztgJcmh8CrPXATgX8JIpi96L8pwkMxCQV65a8deA3qVoSSpk
GUiBtpL5f/uIvcpz+oveV2fvr8U9qrbVRgtQX+Z1SPhZfLtbY9T8NkGCRKxJdLVhWJ6sFXvtVZd3
XQ14DE47qHj/JIcfkBuf1nFkKCX9QKpYHKcDkiQve/+++CzKV2ic6L0zxPzmJrcUu2Mpd2qgMWl7
UO+ch+0ivJDWGRrbix8RS4z+d0OEgaxFfZZ1S+0P9pjbISP2WzOFAt5KBwfMGF5IAHSU6xPSAJwg
iCC1KSKuoQE69EfOh0cQt/02wTY7PI/03kZdRvo4flsf81YnADMshn91GU75MATcluumwwfOez05
z6l1KL5DLFF6DOiRhTt6bh1jDzs3Wa1WeznDEPMpqHbSOHxaWyJbcu46Hgj1E6naGGmVwQMSgc69
5lNhwRQlGC8tfyf9jdeyUVUk6VhYIJfJxXrg3Dg+YCL5gFS0DGD8oDi/m9aVT3maJpyEWW6JQYxn
wTSRgmK/o8X9r1YUuBhT1d/Et+Vrj8lYI0789+pXINE4te2NscF5/AX8rwtOpq41WPK3Kg/H352N
dD5xfQrzkBmDaMikPFYhr/sudMz3lCih/+SHlD0a/rpotgPOIUVJwAHVEBom2Rca9dUZHN9tPr8s
ymxP9xNSpeBOkBnt553qaARQK5gFVIXAEYL8mRKqn5NKqDcBBkK77W/7lmzjibH7+uFq9xIbEPzR
GkGCqdrgQr5FVgdgFbwuvyn6HwPjuIbiD8X3VWN2L5aLA+nEKOpt5fJqqfpEcS7O+17OURugu0MO
LcqOJOHNPfhEvKWN5np+c6G7gFja2XBnnHhSbvyvc0P2uDO67roEtsFgtt5bdAsNCoE5ndYputSo
d6Npo0nideFn8YNhcUAGOZqztJxZxURRgf0GUl84uV4+A2WCYhyJrumMF0oXPZENQ6by0QZmIYBD
pRxZ/m8MFhIVA+yDXZYstvb6Q4HcLPHUz2HGSIghaV6TMKxSHlV3OYNxDWAG6L+HduyEXzRjwxVb
lo46A7JG7iskOqtXuhe8NfxA90GKL0oC4lJcNZkF2RLBb1Ax/HGmugsdu/TCKt/aQQzv4VPZMzB+
EA2o0/qkCB4YoqVoHowvahoi09vLBJooSdez91HVd39tzrYX7JY4Q3/thfT+PvWzmYuF+Jsp558N
pMy/d16wLhCDWbeeKKVEHo7Hz0nAD/FLlzqm0kox/kDbXmzfGe2TaC2KNU1rpxAnye6CUzStKFiD
SMPwNg41fRj0cLbQC1Ac+YyD/IHSegpY9aliFhi9OMETkPJjNMX7Jgzt0nLTBNZ2vjyxF8Dy2UP/
AsolETnC9jqjrD2AL4dZT+U7BLBwfA0fCYJLeaKV1TqWW7yVxariS+ocoIlJZEvJ6Z/DNRXxFlO2
5JNKfM0QMDc3GENArFr8Uf/iUI4JwyoOYSFRlLk3A86rNL7Ew04YB3/nHa2Bh2AzXHfbeQ0VVRca
YhjcFrQl582CfIWymYmwihPADi7LRjRre9yyLDIHNleo2PFfSfo+NSDD4s7YFGNdk5HAwlldDh7J
W4/SQJvA25cF4Or6JGPvin/j0RyBIu9ThJ94qcL0sq22b0UEU37gcMyG0NFy/37u2QK4KnwmLNrV
iEo87VyOLr/EkdpoOVYHrXpHXTI2bmCJzvDheAbPq/032gzkjP/Q+aSLggv4Yp49bsF1z/0Kj8Eg
YrjAU5x7fO4+Js8RytdmD9uOZSfBUtjtGpXOu7wvI+d5Omlpl2WhxtZ9Q7Pk6myeLoQ56zmbBdaG
GrZG6fZQExKH8mtFqmnPtnKMX1zL1V3WfimJRDqG8j4eyXHknNv3HGbV0WsSd9y0PBQaDZKx+9PL
yWGTJea5IwfZoNYnzdFhdlKVRDUvjxYE8+3r8xnM6Lg9dB3oerX4f9mjgj0fwtrq5uXztwjEckEv
h2fUpL9noXksWf4+6I7hzIi5csiaS8Jj4F53pxvayeZQ3f0sMiOFaBcSL7WQHkdLnII8xThOfBC9
tzS8ekHojyFaUzvfNKi7KU0jhbxzmg5NZoGG1hPNPbiyfYVpfHmBeO8LWax3kOO8/zjeUaXDF02Q
KyKTwDcNfvxz8Jla5xz2wclmhqyzMcAuSkjkaUxgbiJCnUEWgQMFDs3zrfBYhvyeLmgp5kuInI/E
i9yxdhGDxAFqf9a8pEVLrsdd+IJ1r9Z3DumbH4dSYUG15jChyHL7DfDi/2VUf/p7zvM8ZhuMj5IP
D3lFGO/oIGW6n1t/irfLLLccO4Vdysc+4VIE1I+QEE+4liggBIk9ZDyVw7X6eR1bNZxM06gL7GmN
9JPxQNNH2CAqoh23VyOgIAlb6DZb2Zl+s/YzWlC19H1jDe2T2Ws6zv+eYcLPqquYKcoo9O0LaLXt
y7WuZgQ593Yhv4c/usCqmgOOPB9wQ+koiu7S7/G0PC7Y3sUTXCcggnPzBIDZKJjbM2GpIrSsSLr+
TktNSOGDYS0gxOTvzPMIvG7kUYDB+mHhGLoUb6ftyiS1W6gLgNyZw/sAsHa1foGncUTyrA85VUek
LlwMUpf/GDAYMiF8mkYifZf4pm9T9YOlNTFykXEuHYumms6l3LA/mzXxjPTh/AU337AEXgSCymmm
NR0kdyhPNZjLWFZkJrjcUQgQ+uhXdTeK04lelmqs2ibo6KwXVMCI0YVpVjmqeIuW8PWlYIse4qjL
K8xmm35NipSrBqs4jm/VDtSvCf3e0C4Z6V1wDvd82YTV6qWB29+OtG+iqOWnGpmBPkAvRxQDkffB
jKe/JJwgoV6XAB9X+9W9cS5Rlc+qQoqkoTMELC77Hkgaeq4qqgVQsh03WCEWhDs7y+6Kjv8ne3v0
KfSHRIY4IXz1b2u/9uo8M23fZmys18Zr6AuzKZd1CSKaav45La/4NJoTWq6GtfDTz42LWOBQmy5I
T3C/yckzfQnberV39RjUw9896UiOptydhymUXJTCP6vcDZNHhWsbr8qsXh1M+SstE3VyDWjWz1mZ
HJSS5qComnl3cYZY3Y66DoC6WtPTc49q+HAXvIRpWXqcTqe2TcIv398amt+XROcekGAhiEWvJ+eu
TXiivxre6Poa2uKb/zh3bKlnDREnZC0iJgromXi5SDENIQdltbtV9AMGmJtHfubEPJalv0JcTIeL
j19xqtotiZ+FGNAMpxuw8ekbRaO+nmu7mfeAzZ2oaDJbgN8wsFY70CHqScCfFrcp8eRHYWPXK8JA
SGiXT0vZVYFdaVEwIYhYzxJCs98Wi/Qf9x6rg7j4e1YTP7V295UvyiYN9V5P31mJVsbwFcoOxt9i
2D5fT/SHqCv2w5OXS3Na4WIx9vpxKVgmr5wEF4kTM2RLmWxzCmXYdqt/eg7Ftqe0jCHjee1zYr/5
hamfWIJaaQVjkibBCbJ1R+mhwj3lwRXXtyZh6/JMbRigHw7Id7kguPwXOYfFE18O8nGew1BA6LeM
7phmRVaBKdZCxme1mtqleBaMKMnBEvrMnUwAUdUhfRZi+26qyDKZEXflgzpfPjB/DKdy4yHT7bRk
M8LfgsvYwRPOzaCeaav3P8YdlYXvMS+5NQYFSUaPh1hmWn7oAAthLjkSUItJXZ/lmJov0gOKSual
aOani2okPZpXSBOCNWaF9SfGMFtxWtmb6tPgUe8dgBrttl2vxdCMhKrUpGODPn8ZIRRHZxhR48O8
sFn502yeoMELpy18jzikXMCx4J7iPCrlpZYOf82b5+Fws0U/Le7GDXlMuUSPu8lfufVM0Pzuxttj
ZBXoT8Bun3E4eIf532rQG+QnEuEDRqK0AIpRMkLcaA9QvEDQbIwz3T7xLAGmbaKFf9zDKldDy63T
uUNXof7499yyjdPZuJ323AOlfICfnxQVq0tVZqqNC3fzOX0a6GZwMV7pZuxuAYVt6smeAd5+Mfkd
Smz+Q2iNT0NpD9Vck9nMQ3UDyUeh2fnC7MvowbHgfX6k3gFDfHAFdtATHvJSIcWLtPOde2FRskej
BH4gYU7idfbSY6bfwDTvRdM+nYlujP2EyD5k/Dygs7G3whu1qjuvm56hAuiJ/LeJA7US5/y7ACYR
rpFUB+hIJqasDHZ+LaKD7fDseKwdiz/p9uczLINKuquLYVtPbiN6tvlubY0kVpno8seXtagY8Cfz
DsKvfFbxmdx6BD54JXGZ3cuFfXoG4naKpvtdSX0CRYXsC3E0CfXVjYcPll3FWH3n0gYm2VAwAkj0
2P0WLX+Lzo734ksJR8OXsRcgvl3iFPZUtJ4s3WMv3Y89d6te8XZX0LzPNBzLrVICrnVndJNsdeoF
IC9fNSRQ2iV14dSWFO9/g1SJsBZV2Pp4bkX5aZG9dIgeEo2VFx1mKTIK5DDjVQfzCkrDXOgMxRAi
6Rx5w2EmXrYaYIQlIjWEAX9I61xzwuwRC0bcankuXW6W0rUi8NGbLtOm7IZoHW7N6pI8iZR8sNYt
t40XSzKp9N8Acx+Kdk3mUTKa4GFEUmDXs4ai29jqO7XgLEVZMiUKpZCIg9stR73lpW10s6d782DL
C4JEjgip5eduojXZn4QP/t7SfIv+NF2ybfY+C3afm2Wk3iWW9V8u/CTXOAumdmc32fTDxu6vjQu3
vZ7DUCQGNF/Oq+cNe66wFFnIDQBy2N8gK0gP3CHkaXY2iF8bP77kzK3pMB2PCdxh0/2zVG0mYt6m
v/W51a+FVxeb1IA6+SxhsIVMhPBafaloS2AHSbvLaM8DC0RSEqyKtbexQwKq93Qr7zC79FOnwjpW
bRUb46ELfR/jRRIWDosfG4A8jhfbvN1NHcBtEF31aI90I4OTxV6hRWsn2Vio9nQOswiL6XZNMGnz
v7eTCYnf8CCJTEyPSXH7HrJvOByxFBWq61n7t/uQEthqYZu5K5duwOjWhtyvllkWGd2AzsFeA/Fd
ySrm0Usnd0NolkBJzHm1LCNBmZsdGwygpj/nDonlLePDZzOglaYsQzIXdPX9lhM2ZQ9BdOeDpdiR
OS7yN9WyiwNaWmTltrV2zIcscB5BHf6U0qpfWC2NvKSiZ5ZXVMDwxQV93bzoVWG8CE3WXcMYYqYU
PoxJiO+rDKZgNU1S0+KFa+5oZ7w7Lutfxnxo1ASLBUv+DIHcqpIB3CGJcr8YiYoeX2bEsosTYcOP
IR6orZ9pICYHKcXlTXeQrYoLDpXIcU7+ZL9zHJHlLBIw+fdQN0M6qZE+5DKhiExWD4Mibj02Scat
S2E2nJy8R47Bb3z3ZHwWFCoZG4zUvY9AdHhnwZF9rXKbEVK+mOPRTZrDmRrjDx5UMXeMEF0UTFQr
dtI+Skg69rIHOoNN+eBl/IX1HfWXZSJNkFnSs99YuPpW+PlMBpO7aSBzyFaS8Zyx5+HR+OOtVuqB
F/Wr1ht8KC2k3jgF/q0Uz662PThFWmRQAkyWTh7Hk5pVuSjxKhBbb9OHwUqu73uSpOlR1AoU/RrG
PUKbhVQ2kKdS+k5PZvKCxBqdPCX/YGE4uci+YYYjCJk2C6Jf8OYAd56Ob4RcIVZmsIYOZQ2wPE6d
BVgoGZNjn1/I6qgm1SjipCXUSLKvohB52b+qBEjorBSXWsnqxsLuihgE94fCg3j8BjQGaWe6UNI+
zpyIf0zhVlU/hwopfs4cLhZdkMQYS7Hhh09zUCIFuhkwQf1KqyKy1GOT2SZ/7V4nRWs8yqiIKJLb
Rq3jlLIhlktsYwDVhpxqlLxr2Z2+au59NPEOFLwRBg2yKW6EcV4nMg2wgn3lbFYiiSJ/K43pAoNf
J4F2LnVGkkZmVCRhu70yyHABtsjo51Hi7dzOd3wwyH+D1+rP3HI0Giqv5lT1W5/87ogrMb/Pu4vo
yl7JiEoCHO/ZZYf7+FVMmHlz/QHs60j+JfDIiF/A36IAHZ5x8aHBZV8zdc7RxDJIdcQ6FHlhSr6A
y+gubqRZBtfCgqeUQa8VXdkQ9T4avwIltxzfKxMHD8kmHSmJ1mMSCDrxE6AdBl1X6Wtm/YJ6xDNt
vl7x1hhbUfcuyG010X7nLbraTygPQf/QFJG8lcDx5onXs/1GxUAZthJANmx87rS3zbkEJtyzRYbc
j1SGIzxgw2jt2uQX0c2ctFWno0CHDrslFx/fP1gTO7dR1UI6YpFTtv0v1N75BZnUm6IHIkMrKOP8
x/Ic9fqLgYkzQIH5wC7GU8euZ9Sv79DmoE/0+xAg+x9jcWDRdt3/r/LXiShKBW8UnaC5k8eaGemp
Kh/KAnlmVyGgkcWSYy5xqIb6akMUqjSzj5WuoetIksat7FnNIJHU177PKLsfTzcJRQb+cZrYy9UO
G7Z7qvLJCBkaWlL09W1SKzSfg5AJFisaw/ClTSX19jz88eYpNGzT705Gf+dUOEjkSisjx/h//BlV
7uqTmmeNwfo2i88J3/mtIgmZEycpBzrwfhbFQcHbSU9qPdwi07K6F4/dbBYomkkjDwpBRviHQswq
wkNNctle/vtEnoyWB6Jmpain/kNwrqFfmSg6Y/ZfMzvN2D4pNPHTMi5/6LcdZdaLnyWjbFub2tjc
YCZo7qwCYO+8mOAxt5v0zFP067dCxmyTpq/qHNAOMXXaCEQpVLE8DhqDgZlaPyNpylJy+SIp/3qU
3LUChvzFvCm/XTidAeUW+TW/mdIFyBlzsN8v6omyunhprbMusEftxVC8wEOwSyeLbwpmc+eV8GVx
EBUW+6kHfGnccqoI8tSdYIYFn/PC6vk/tbJEGi0vYF7EXtrFV/HqxKfSCHqu1mgemDiowDl5g+g7
7oEGCkA3iV9Mh6714i+3iXodlmuHi9rLI4V76CjL969mO2jon3ny2z9VGlWOPKadgeNbF8uYrrri
UV7PSEt1k7GC5SjD7bIjVMFOi0H6g88LOTu31NQAugtRX9rEs/BuZ6BsFRVWe1r6SAseHz+hV662
Xw66BH/Sn0ukzHtsNr3QZ2z/wvcrsBegidoryFRGzYb1C5qU9tfDiEWRgqFLnMd1MuUjiFlqf4Ne
BcG80NQ4pWW5nCTvwS2H5633Fnb3Lsuidb5Qwa3aQFshQGKPx4KCBgV9izaJEfEppcKoVWE85Z6A
06PJOD1DhMJGsE8ORGDQPoU9PN87wjJO7vqssyo7akZ55UXsx5CUkVgfpcoktRTTX208WoiuXQSb
8453tSu8G/oeaYhtFG9giuyxtMQCPep+AZMxvmZ8raMeBPZPa73vAt2DQKvlJAP6TMdDRSfqFhrT
u5wOnkMm6jZk6xbcHbjQxrqk+eDHgyW3mPZoJMLHmZcWdvr1FZnm7cNtG+Sv5f0G2OxVaZ8/JcbY
16B/k/gMwXkHIUIH+KG7RukCeRRYyRsjKsZLRjW6iZkw5XvTs2ZQXpsJIxbjYUr7GhVgsXBFUOFW
FKSmYO/pcWULZWVoa4GLaBdHTbZjC4DLjHnWgq/q6q2GV6+z8WMkn3TuQHArEDSEF/5QSCbHr8Oq
hMmC7koWlKfEodc5TwQO0OJwpgPP8hhUtE8nbaQaJ8LYv0ygm02Y6S3IxXkohSBR37zkjf7P3iLc
kG41KEdhqsEZxSIUygysmZfpPGzo/s2HaplfZ3DebokYfRTcfGEjbKBx4C6/NQO7JaJsnY4/PeEj
viPJQwVjAuhDVUwTMwbJbfyZov/F0dpnHrNwOC/6LVaeh6101/uA4dd+lKq/Z/VUWZDQlGiQ3Cpp
vGotcd90tHQ/J0Yqqop7eDYYy39la/jWSDq+ucYvHXzbQq5WQKViIHtD8GaurWkT/T8k23wwbOQN
e06wXvbIqBwZgloFlMfLfh4eTAjudulrRh90RV7JvAiUDXqzidV6pR/Q754GL0F4SbTclHvOikaT
88XbrHFbmqMfHd8RFAxmEKzQak1vHCsCxkzBDGBAZ+33IykOsmiflr9xYaQOalpRRKX5jPGZiV9K
1y97l6n8eSY7nC4v7ZM1prRt26t79pIY7wKYcVImxGiYJ945Hw+zlsK3BcIwbpCLuDw9y9QNKNwL
lxBvFpbYQckpaadN+JpSSrQG9DT/1wNUfkUuLrMsdT0NTOzWDUBlOo0QzP/vAC8Prcdz0c3X9XQj
MKTrIxWmHtT8UMJjg3I6Fiepyn6yXLeJfiqsS1R5c2bjXgY3mEThqKejyj6b+amcqojE6cvq0fAz
oZOaVZZuSlVc3CCU/8IIZVeH5AAN5vWJz/D86HAxDFLzdxCtH/lUaI+8jLvM4QtC6NzXxbWM0a4W
BuFivbeRFTiexNh93e+RPn3ITvdEjkyuSGtCujwvdF19d6PZpCWPnHlhHY4jIc1kwg2g5Ms92D63
/QAsuRiEjBnSAgduA/uLrAHKDsN0Z/iNL11eUR+HosimXMKePTyf5Qp6gFkEApK694aYlT0E2z5Q
DLrCwtEnkX5PLQeyyys1zIG4t5AjT2E8FLCCABfZUJNK5erzAGtdE88EYB1MNrG+y+cpiq8I1hnO
S3jyilfvLFtCpbg3y9XiVECASE/HOEbbXlQfWJaYBUhYLB5Mh8Rr2GdYGu/Yn3hPMPJPewDBfs/A
MDWoKA1dMcoPnfKxSZT91Z+uFEccbeouvTjYICL/y1sZNHQ2QC4w2TNPUF6KvgsrnstQlOvdffCc
o6Zi/QY0kLAy9j9PQ1RgY2xBfn6X/adu+89IZsJMgusJ3Qd9ZXsUNsZO+w348V5N7lp30iKriGEb
+cIGfHRM9hVfn+yHuH4NYtn99YeMpZZJbnBJjPorK8u7l9rMlSRx9yLBGK06AeZCWaWEUk7Wj6h4
L7O7tFiHC+6n8FlOyph0GRn10vlLAPW9XEok5Xlm7Gx4GT+dutIT6URHNMla8h9yTlBa7CLD4TRu
5pLUTRdhy9UWkjEYU3zy70gQkNVPh5ePep9K20GtajFFrifhcXPJTPRngsWqQX+uf/pIqtVgi5nf
TiE2b9B48JqU50JInDaGwLk0TmLJwXA81NAWNtpZIBi1P9iCuw/v/ufKKzl58oUqmf+X2uCtugvB
i0gtu41vJwPMXBVkNWWdtifiaYG1fF44gNjcZR0yKpl5Eyd2UL/S6UcNP6zS1wyNES3YQK7iZXCK
l0blTQULul+GKqEEfLd5RgOtXr1k9l80Ev91Auv/fx+K8ySVrGlWQWgoX1TRsoQ5Zv5xswW/64Od
5MTjwG6q8psfa1L8enoISw5jLHu+BRnT7uQAZ+5yMhFX/Gytgv1N3GneApkf6glYh2BA4/eC5W37
RNMubaLqVc6FbyJgwjrezmzkDlABVlDEVLgcb8XEfTUVucH1tnhlTstqDkIEJafXNryQq5kNCMdA
8fRhZJtRvJsyTvw5xEhcTbfKMRbigT59KS5bMbedJjtFlZYcSeVcmz6+0dhO++h5t6kjByjtlN1X
HU9D7SGIfSsN99YdOq1t1oRqffg8WP/mxmGVoTIhtRe98otjYfTfXatp3uI4sLedcFsNbc8qWQmu
wTPG4pZ580yNMgw5x/1tmf7H6yfsIM1nDf524ZMu19yzEn4faEEypB/fn3HDDvrIAEYpOkkKTnDd
Z/RnaZt56OZNJDUThBbIyL3ZuNXPjNDDApjYimP5ajlX78Ifk8qVhVu8GGmmhpZKqJX5x0OK9yTa
lKFU1p1tMrBXnIZw7C9cpEc39e17XVXlV9QKMfSzraFEm5jLb9mIy8+pDMyUnfiqiJY1duHpGvnG
OxC8/P7c5HOkJpjte9DRCzwGR4rLzQtOEGEraku68Ti2rCtl4IVCaRsR9isYtKZTKd5YInXCnsOI
ZYCpStL2uNnfeXCCmbVFuqYIuLRFt9Sw4tDKbZTLNWsLoo1x1H275nNFwV0n070jVWgRbSUS5W7D
kVNfEcSeGbjWa/RZl8wGx4WEdgRtzUevE/Os2DdCa/Nf8mypZt+m8zsxz/RsxOnnP9f+B3tFdQ9t
2waNxkFhwRsyOrN7Rynlg5MMp5RyPZXUWMiauBHGJNaHtLDrzQp2y3l8mCs36XIUeac2bk5iEMlk
alVxuabrm+7sVuTRnyK/FOjCfCZ/Qp06TZ/bg/wfNQEjdqWmtP0g6d/xcI+AVSJtn1IjCXWW+VCS
0373ICaqY3gTt+XRN+hQKCDriD6gQzY92ZYeqPvw/S0+4Sxs9wQ9iEevzjf7nwv/ZfSLq2aYqRc5
OUxBHW3c7drP/awVv+tzDa/HFkeaorH/OWgmBdLIY/WX0oG1MzowbZZYbMDH93jd1i8Ba6KlHNqa
jx4abzID4ap5ONhv+x0C1GtGnmwFMYni6EcvY7u/6XCg4HpEwc3sZQIA3hK/Wu7J4WIVQBpVn6Xb
fjeqXP50fduurg0R/tr+MNk3dW7Eym9CLfxJCrwhdiTAv1xy2luyAob/5PDknDJ3rltHHL2QhNJ1
1mDDBfN5HUgHMOt7EC7U4QG9ej50qQGEQDy0mGtuN9VKDkqKu7OaHvDCNsLKoEWKL91FxtwZIPCs
EGXe1PZ+oda8fIs/Cd7oJ8pvg5fgihtDkffGtcQ2kp+/zyg8/i2o3Zk1mWMSgpt7tY/x331x24uU
cid57VsN8Yvu/GeO8cFj/oe6GpIJmACVz3elJZv0IM6GtbOEVBMojsLvpiOYE7OT0v9Lwb1bHQ8s
bqAU3QyCaQ0w1I0YXanKXUcwyL6ne4jZW7AtRjo6Tpyqljdso1NG3LFBp4s0sMuWD8IXFczvfKjr
5LMtxsKwNdmx1j8UvJ4Pnscwt7z49i1M2xZ5yG4yzPV8auA0/1M55l6vg7xL55Zek/xyGENn/xOA
4TmWV4CsW5FF4k+tmldG4HnpZyLZ8y5du9VPJFSz6alF7iux90NzZEHqIrOau/IAMa2u0ZEjY7G/
CTLeQYE0+djdzje8XLJDX29XxcGUjG6CZSCkcSrnddndhzboAjw9HvKxv5vkwN56DHT1qEXETv2m
OF6usQ8FY82PnChia611+i+d/tKI0htH7iWcdUne4yi4B1PoypY5dnMxnEp976fDyn9ivT2uedqh
HyRV1nOmD1vZcoCiBLldW/ICzHjXw9bCcFQoZnQFUDDyoVAVoiwLs6KuE3skETmg9wyt7IxXaE59
ujgVe+ECsKj3CjwNX8iwdIj8pNMFI2ykUTzUZAFSu62V06iKs0olQeRDvVcPNsBgcFBzwvs56da5
wkR2hnVrj3knPwPLQ/NFfyCwqcz87CPLblVdrNyL3vRvrXMKt9qwgbz9iP37R+kFuZXPIQ0FvrG8
l2RBvvoSv17hY1hO6NyPtRM6kQ3hHoCPJqVw1EogtoTjnb2uNuxhoqWo7U6c2/tU6NFUwFQSacMX
cr7QKp4GL477fNNU9wq3EZK1gVGiDRVnEjtoL0LXl6Sfuy2u6Ye0re49Kt/nOd7rK7WZn01fESIt
geiQPiuq9bOwByXaO5n/9KBawNTVddlnSIiOeapTSrj6YFTWGEHHpRWDf9b/Zndlab9yXiYKjQ+o
4lrZsJUEnMwxhGl0enn+SQYKBRyjtaZiJzGV8kHh1J6nH+drlMXtp9XOr/FDkzAq4ObJPg7VheXJ
7J9vG3zvuhNTnCRClvEaqdzCwir/kf2MxdcPvetPfw15ZBbPO5gDawjFbood4SBpC5PQOfHjnb+B
WrLXo1VfhO2rpyn3aWTNgMbMu+UVFJwUmYMoFTF7aGVNf61YNYaHeIYCK4Wz9WSspWNCPCGkhX+W
HMzJpJeqBEm1QF3MKCVH+bZo7ppQxMBxRVZzHQUu5aMbvGIKLAgzk883jwAY7a5HqD7hnAEzO5t1
jGxZwGEjvq8HStBpCkZtAC3Tqa+xtAbgFjAZFY31LAXQXg/KiBQBdtSocrbYVWy7md14kV/GA9nM
JJwBE2ET/JSrfd2lEPlfawg1t5+CHebiuRRN9VzuXD4ZXRaCRn2S2LQMoVFBJ4feVODu9hJB91Tv
mSQOAcQ3GG/3vAoNgXbv6vQ4DQomym2TQIQz8SUfPVZutfWOlE0Vd3SoXdErERCuGMTR2h2GnqQe
aV0jx4AtlDzwlnpdYBHccrZDZUY9VWjIE4m9wELwbw4riOmVAyPRlxUwC7SRzp8YA95HTD3Yy0CF
fCl4Qqxj+3BnazGYStnBPnRlsoMrmLKXRsnfZLbi6hPSVTwHeWScWKunHa+6jLverb6JRNdrnMTD
4QeKk19AF8ZACR2p47XYKftmA7+Qk5JScyc7g8gaFx6XPBJhmMVfhW8qJhLlcD0vDiH5e929qylR
fMo76kzwok9lnS3ZJZg+5C+iBkLUVWqmdN6YVmEqAWGV99T/5mahvZofq8wHZPpKv8w1XKRvjqf6
NRg6wODPWzALKEhzwj9aE+1A9JNvkRtC+srx1YHh0/Pzgi03GUE9MyGRlZ3/rdqXSrGX9ymY5XTG
/K1E/6/lWrofPWHTvjXOoeEMZ1NQhCKPhzodiqkcjmbnTm96jKbw/v1eGzsI4au167/SM8T3q+Jh
fnIXIxzOcpIOBfq319O4ssOkxys9ydq/Lj+HrzFFsV1RThhANzfytKjam5I8bgaf1q7491ZPkWRG
M0ikPtFJ+ic=
`pragma protect end_protected
