// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HGA7cKvYtkMN8FCyKoizurKt3vdfdWHXgKIDHiP2u4PwDwzxffuunl+XE5bNlCwx
kAL6msKtK/oTkMd+DGkUA8KOZg1aScLupGccAGUangto4k0NewrBoBvk2o0GLCwU
fWotT3QxA8gXBxDjwTJDmYbg8Fc15Tf+GOGn0kRxW5s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11808)
HACpy6H0BPaDz6rSIqteZ4aoDQoFPQ2i+6QRvI1nYa648cDL6Z5nCZHKKs+V2GrP
xg/iivz+ZjAwRzKrS272DXFRRvdiUdrMToX/H/wUpfhhvjPl6P0EbnnTXogKaVQe
DmmlnRUMiAE2BidijRNo0galW0tP32tV3Gu0GqPTxJM/Ndkjpkbubvx0OhWqFmuq
3y3TZUA4O3pZ0beZ4x8UmEmnArpcrzd3Su79YbdbPtqp+gqbnbQOXmqWLfWFtia6
NMjnCFhIWpRh0UKJY/TYNO0xlgF3Zf5juDHsKrVWziXEeQiH0HKOInWK0V9qdVyQ
qID3t4o68/wJrBI0IJ9rxf3VG1ZS3eaSSrO3yIGvdUPU9sJ9reaFLk0cr/HSiGMp
DXjoWHE9jxSv6LIZCmRssp3DGXzH1TpA/uXarUYGi/MgNMLjhDHCS+cavgWRTgkZ
wqgiOlQvpA7zkpbrmYwtMm1Aoo5N34M6TGt3h9gg4lQjUCQaFbXOfydwu0k211cf
OQnEE/dMqMlqQz3K0z/jmb11KLbVxDGqvCxiD4zAqfap1dqapaxOYXOf+FoWfu58
/MoZ6UGvaZ5BX4cjuK8+RKKY9MCyWb/7prNhaSqCx3q5E8otUuP66HVTayn1xwJF
it7JtZD4Y9BlUtX6lTbngAnwfVEvdYkrKS3L/khD1oasGsLHKkWafhTqn0t1xvxm
ExXEWQZDeeYegRbNSguTcsWEfjCyxge8+UZYJA1QQYjCyQc9SkTsH7x4WEPitIyR
i2vSt9HxYeajMzDG6k8yGUvx0i84nA9OUnudYEeFvrGvyXHnJbNv8Vsdfck7U2jn
orqvfphi8m65mupyTXid2Gsw/yC+OzgGr84TIgQN4v+rnErR5mgXIpb7ttFkgEfV
FEJro3i+6f8sGXO9gV1Lz4bAxlkajRZB4aqw5p2tL7gle59JciS3yi5SdBo0xtP8
1wQCsJHmzuK/MYx7yvrKWrQntx/WWAdyFGMXCfU2003PWG2UYZVFIixzPeHhMRzr
f8vI2QBRdJQvM3HS8Zc3y04vRdkXLq4hujZSMM6RnCly2jLXGjro8j4Zh1fOk6T+
zH5qzBmWDT/gez5EfUNAVc1uaBvtvcVUvFF7li1jArw6BnF9YYmMgRfQUKd3ZN6p
Rjn3pmc4vuap30SY2CcvvH4oDWVBcf0VaDbzhmo969MitDVwzPOwfcafBzUbf8B0
XVJNaTx2UMm0tKiomkxBk53QSzKURtztOA5LCBBTUTspivPK2yth9KgsIU0rlTcE
WBccwGMdY66PMShwd0l4ttXtKmarhVvGShuwaUNGaGLWe9QD8AcETa1qcC6n2ugV
mKjOTMlmy7TPNlR5MVUUmRcH0PQLvRFGA7atxNokJjWSkIHTgcakOdA6T0a9HouW
C/MsvnswW+38nbPZ4GkkuXTPuaSrLNx0DclsdktdajFCBd66g5I8VDwAjGwCh3c8
V1A9qrKejvgcwXFXRl7Z+bGTXBWArP9T6oX9Uj/RNVJswmGqgk60PFBwwDh7e6TI
0YioetwCYQHZTgs8buk7KcU9jt64BOP06aUJimjRqUqDmcz+PgJC9JxFDYuDr4XU
dw97kYOSHcb//jIYgxQEne7+KabBPBYsIvBl4dHDpRIXoWIFGF//iC3KxlMPigJw
0uC1+XEsvR73IJObqDD9D3XLjtRqoC2SbPg1eEcekNlFHtZ6Hqu8r6vti+d0Kfki
K0rD9U466qJzaZSlnmkeWGMnpHcAAvrx1QOIQyJF8kZTdR/V9KzjJEhxROBd0/ez
q78Xfza3w6R7kTMt+muI58IuIGFARRKdNwTGemOXpBhGrmCuRJ58OYpuc7+lv/st
oThGuaYqMP0urS8/BtokiKxY+9K//+C2kay3oVSA+ETGVx7dEPWC/QGSZ5/BYArc
JimgeUkEO2CPM6FJYKgtrTlCLZyiFgrpPI5tIKmgR9VVdXvGdvldMcIiLXmwUqFk
zspoUQfZgXIXNXPCnVwyUQiEifmllalSOGXfnYEk4fbQW4Ho/FwCLES1W236Hh/C
3oYBO1q6TNQx8icewdbo+srKUIyhHEb2rOSxbY7/6569BpeU2OLDEeGlrP6QQCgG
pp3W3Sf0S+3G//yCSiypdznn8bW8rsFsnS9/pgpnswpeQi12NABc7pNWw4tVxF/w
8Q9xwiS2Nf63+Yerplh+fbsuoUVfcbr/l2guo8aQ/xAGPJYTpBn5Ms/ayTlGDa5D
wTFcUVWy1ZoFql9vkUjOoL6d+6cxZ+Tic/0ckITqrQleubQ8Z/LEsg5LuDBmvYMS
DndJmm1TiNplk6RSMdCrAa3bQAiLGgMoWBARc2TwU6LlDCoaZAVDnLE9apHMNZ6M
WTLt3n5MnN6TWOr1zfDrxxNUfiAe/ssxFbxPog8lJiywFGwWDPw5WtSSHXh0OkUg
xDWcnRQkRZYoyKhuVbcp5EU+EdDREbVQuM41iOVSjO8kKeEIVtacz9/WnI0nxEpH
sh5tc1Ea5ebVOySQY9SuETQfiyoOkTNg1Fyrdc/EWCxrxanVtOnrz4N0sjrR42Eo
YEpMyU0aaZmLAOK11cgPLSptPumYPxHUmHPyz/DAW3UVl4+TY3WZubajBCWcYaup
qsslfz5vPAbHVTrrJYsW/VrIEpD8neG9D0Jb33vYQ34Cl6FbC34tnuT2T/ODXdo3
MYrF0QHvfvHkBRBDaKccD6HALeaBR2lgGrp7xqeBix+4HvU1mTwiJf3w3W4wHBzu
HdiazwlHqfXRBobXISREPNoyuEzuIg8L5PNG9ZI7eVhEaYIIGBcG6ug5lrcrWet7
ftqQEmsUW4yz4LmHdqp950Kxoc5qZPmx6qUdT4DbtFTUGo9OPMEDXzV4wyudaoD0
jcQIRXiO4y5kyIlGjs97Eg9pCXfs3vcR2OjFVrufppcT7CAHpLaLOO+7uP7/Rnzr
N09JBRAbB0P6Z6+KC3YI8QIIEWcJMUzUIxoDhOgMjIjB1xISg6bwOXM/TrTw2xJW
y3ClCCNyuSzzjpA+3C2wAtLhZqKfqvTPBxJk1bezNRioVSGXjuH3aXnDUjPHwraq
nsb9p5Wzf5vPaDJGQp2dV4namwiigXDK+GU6zv/z66Sw657QHBwBPRVhFQKkajNz
dMdZ+rFenFtzKqawr/H/jKNdmSmdQq1THCZzA6c18mXuXEC0DvQIeDvRCmLqEKMF
Hi1vpu17aoYFuTTy4oiSxzGGy+1ZHilQK7QllYAucne4iRlYIqB3tglBN2kJlZYA
y1tx3iJskw5kA0BajUOQ9y1dADDk4BiOeyJO9uCog27XgH+mwjhDbVY7KFMIykWl
U0rU78gybIPvTvC8Y52ro9xQKsHDly/k1QXBi9RqWwZcsLQMWr+MGKZjxNUhDiph
2ISvFbY85mT8YKaIMaKmoYDuqkadylZzVGqSfAveG5k6Z5pxQqGvG6RtMuErRW9W
9QERXp/wMHv37eIJH3ISXXz8eJoHSIizbHyU70kMCtfMTVNPehq4T3pl/RD0wbei
K7g2duOheQg5NtQWv9YIxNGvXzGE74v7WUEB+CkpP2u+LFVbzIZLkyWxzjCHLLJq
qt9jsYmxBo0m6TQsHLLbFwLxKzvwiXxBouUGAckxtB+kEiZKKhAlzVdvaCuEn3Cf
MTUMy5yY3ZJkUYS3R9PgLN7IIk/uhRdPzka5l+Y1EjMPtos+zlOUuhnc+sYa7rzT
8moT0GIPbvHnMUaUI63HtBCbYFh1GQ2iO50UUOceOGpSVdMUmnIz9iGfnHqwRGdA
hGm/qaifdKhTl5Q4cMDhv80OiXAvlaUCiPBMcwXQx4QlhjI1kLLXb28D/uzih3xn
6YiZGOy+QFDGEo3CKDiXzmqJMKunLCkIuujxuavs+lajYaupsjdz2bS1L+WUwAhO
r2i8yEV0Oy5fxxqSA+wFMeysVCQC8cfI1Lcdi96j5E+WBFbX4Xij7Zn6zFouO0Je
Ul2n4o9iJs+jc0XwyRgsm2g4/mK36iIoiV83tvxYtKVtBbOHiL2TmvhW+NA1CtWx
YQtlml60odaGVHUY5B+CPqn11T7aWBT2oTy+S0FNvv+KpYREhyEhdNh7fJoiWYwS
vMo98xPBgYQ7lLMi0pFQ+FqpjjUgDD+i8ujSX6YoIOb6aIVP8UocDhKTxY6pJ9/U
BNv9lEagAxIQPkOB6uWEJE3wdv4U2sSU13qjhRbA1/K8YP/tDtuYuWwGKP7yNVm/
e40bZQH3o9A8on7KT/iBRXsjAazYUqzPCoyvYqwlxtqIf/V836fKrGcbUhs+tEZC
sTwP+6a+aivgumSaanLpk7QZWEUyYARLfIumf+oelEWCSXFU8fi3C52IezzoVBGy
KZuwrMQhaH+S7R9CxuZqacpbODQkLBxDO4KjO8KNYpibs+juYY+K60ViA8uPfGYV
J8CkVHSvmI8Y+9lhM+zbuawlGiXQFioPtEtxsbhsSQy9D/OrMVqiEEk9pwXn6KIq
xzTn7sVwQDySbhvuF81hauQT/8pnPHsiPhh9gNI3qHhqoqb3Ppknz+KMouF9u4U/
3/pcKtG11t3V0XWMUOb733MfpryhKk5BtCewCaVe5/QROYLl3NlpI4K3nr8U8Crp
p4YHTgqOrf5FjEf/Ac7EhlzF8lYVxSn1nZ+cc8dTo9tjorvwdBRBSanrWNBrGUjg
gaZyfpznLlnBmP16d+OtF+r1q/VVWg7KYARp5/pSo8dQWPrO90iewVdtsk0GjN+p
ijvU/SzVL+QR+XRNg6o8Kg+v0u9fe2rDX6BwVzskqMvexLpeptXepy5oJHgq1LNh
2bV0gauRs/2PC815LYff95URdsz341heA1ZejWOq518WrQG5ZmU5xEnyBSOVjkdi
5hK1ZcVScyLSDdQMBqLm610wRoyqswb7w3o6OESSFBGfsWEq1KraSFwa/0e81p/p
iUm6mqgp7fa3pBUVWERW2C9zWQ5oIjKEyPoTxcoVsEU01fcA2+9e6zlracC8dJ7E
CVr3SiSWg6V5n+GUUFV5ZZW2bZacj1jQLLUNCGLeYlcJKvCCYogplkXhZ8B6qsSp
3rstQpADKurnkGhRbj4t1hhRP2tFmfjx1/fg+tq1BtNzFQhAHY+ms6IMxMTpnXxa
BBrDXpiDYzqvyLTxR7DFShm1SSNOgwwYZ0ocQ2EWirNAMOMZONWpMtfY6oyvyXBK
vnvzf5DCYAULB/4RIoohCCmmhku+O2QUR3gb6OJMC5YCcOMNoDMsw+5lRXATpLvl
I7uzJ587aRL8fDxQE6XKfLVv+Rc5pCAxT9EV6N045dPBI2FKoAh7ejGzRdpVcxEL
D68Q8tR7Yr2tniQSrdEsYI6MqrcIt0rhj8Q4J5am982TkZC/nGSWg/aXIi9rb4k3
KO87rRWwf6UfKU8mlbVlCvAYXZ5MvIUyH2tijFQJuQahQXEVfW33iEhdxY5jkeuB
qiCYvL9SaW4Sed1p87Z4tNOk6GUDLo14VMmioFZQi8ZuN/45D/dwKKv3eLMH5BDR
2jXZ13IFE6h5L89o3Yld1hfgJIOGe7m+cWVHeFS4qSKIYS8XZeUCXTiPMljp+dpr
9PXezIlxTDiGx+n1O+QfDfk9eKC7Oi5yS1qEdcE3XaqSmS+LncEp+ozklFWV7IWt
nAtAlOCBPz4MOzLJbmPxoMEzvfhIi8p0mEHSDFxs9tQotSVwg64Q8F048xYFuQp9
QhHH6AmpZKQk5JfCXbTMYUN5bKzi9toxXvUW9yhqfL9dlwFgXCO29EoJJTpGxPO5
3YaPIyrNQAnFGFthI7mFxsPW7x4DcYeN/d/0xtvRqriVHDCZVpWak5S0qwpBX/c+
QSnIbwTXlfNzJObQfzf1KCrUjdxgup06jEF7nllIxXPz9JmA1httXptP36L9FTRP
SC1+kvY6BKjVEqzVYGGs2kwSVygDMJjLImUrpWYU3kEpZpof4ox7BCTK/1Di9e5z
Ex73tucBQY1HJlfgNnc8WR8z6/KLu0u2Ofi3Jnpvif7DXRMSbDcmPogFxtqnrgrw
OLSEpUPXmT8bt79n2Nas7//UTmEvrKaRC2OsMc1WnLNo9lVcgqYiSID2yPMEkadP
pcTEPhZ+LeYjEJV7ZxDPjBxVyQ/4aUDk5Z5hEi+JNOtzDYtq10aLZRTZOjwq3MQn
olYzy+YL1yFAmoPD9c3Qk5yzg8LBSnAeC4sCwKnzCWikZyf7tnkgi8AVR+tAxDkW
3j69zZily66nmFZp0SMYd6xrdqXdukM6Y9VHULrvAa8I1rKdHOFoK71y1lxlE9Lj
qHSF3BD5QbRm63Xl2zsZYBnGL/4k7U0oOloq3PyHTUNk2n9qTB79VmBbqFbYTPKm
x7IWvE7XxvSV9nIM6jfjhK9NheExnE9jp0uJUUBge5fm1q6eeO/y8Z1rlUFFNbW/
NR5TG64kJMjZ2zv3Nls6XFUvxH8OXa8ogYACzHeylXZFU/jP/iSvuSyOlLNA0GLl
9CsaBkSp7TPD3al4PJ/7OUiewomNTEpHEQLaJsW2LlhSSApS9K8/Z61o+o1rQ3qm
rGv9utGGY7llino0M+uBflJqYLDzCvfr4ynwy6nJgySv3346Jniqwf977QEXOzcl
ioTR5Vrb+eNgKKRXGyyWUQ25lK6ggkyQCaVBN66vikylXNG7JLYIYeTLFUHcE3Z8
/LOecQywsN2q1sFNX38dxz8sCqQk8ivrfZTS8tZvEWYXil35iB6cRx6JNmK+skQu
GAP4NTKniKAZHki2ah78C3kHQUmerXHzgUDQM/8GueVjzAChN3uZpZOem7JzW50S
/E8u4V3h62Dpi/XR1TGfbYly+T2gd//zzyhvE6yGiAi5V7Qfyurkr6wpMnYpFwsm
XFLzJgLE/8Dz70wIdG8X3+fpqhynQfzRlhKzPQ6J8XUOkSXueMKGucHUe7mly21g
cD3+zSOnjJA0+Cjo029JW+2N8F7J1Jf+VRSz7X6IyYJaJuoG3eTo8EgFh5pmMgCH
+yg397JQJM1gaJy2EHCbqumyI4wZS3rO1r8O5EHve3zAknGMG0nTia4PMBmmxRna
ITo4Al/XFjnwgHI04TRnlg4kSKmIpvW+xDWop+ousGLO1OjlSonq3X7/FcJkBz9S
U/JDvB6Jz9m3k93yWuh/oqPD/hH//HcQ3IzYkRiSksAPt9BmHNkcE7XKMTgqRH5C
Xhn1K0LusrZ+dXL0wGfrf31dq23VHU/hNAbvr00Torsut8bLS8+9sYW+eJUKzInk
3PUMAnhJk7mAxRdEdZt8+GGtCEdU3UGS9OqfaIL0wiZVFnxMM6vhye/Z20d4HGP6
rwPFsERurQnYcqWRYmKILBKzWhED2Dv1AAJUmEl7Cc6dbmbZBLM1kezWwxdYC0rk
9bIeZD9dNRdHNo3FSRYTTh8UguZCmakt9eDNcYUx8ESlnuqOtHZly6RjmMyaX1cH
cICa27s2zr8ad/drGkig4dTForI9Q/R2uqrcR7LwbmnIr7K78tyZ9B+sRoi4+Zmg
IGSBI5n68a2o6HJZCqIPwNWJXF/ZReFm+p0Jv259SpfyqTNogcJ4K87VrcEwMT/R
aW5EffQk9g254gBfwpYd8HFGe+iZe03gYubyh/3Qw9YFGLdmyGXc6qpqphcB5qbG
+H0QeeI8dZ4isjYevHKJOPk53HSSoC/nba8y9ZdOmzPSp5WwOrcYL9mAadNlXH3+
uq+MEocdDxN/Nuj0IsT33Cigg+ksmUlL49OvVc2/RMUSAZIZSwt2vTcanjM/9xG1
uMnx8+/NiZFPHZ3yV+rqfgQQkXpdmGjAPh+mBBzcmUvg2wjahxCLsjgDLX1g/6QA
OLU+jfUpaM57ztpz+REtKcGyvTjPmCWN6vUXi1KbSTBqP+t2R56bCziTjVkQI+7X
viMzaeUyRj3dJTFA0OhXlql7dy7RxB7RbHaC1MKYe4QDa6Awv13piIJbaLU5r86h
Wtgqz4/R+3Y4lTt5ZTjJSPtvi67yZoCabiufnqIajkDvKQ8q39/f9TWu1Y4iTd4f
NbPYkonPKtJM2J6oTQc5wRZarqwEoP7/txJQHsPB//QhvjHGiThzc7BPJm6XjX7A
RifMWqLgG7T5gzrg9BtmFNupRQd16686tfMMLg99VIWsH6JhJeHllfKfBf32Wm6C
Nz6wkNh1AAz/v0eoo28Wu95xnt0cIzde/3Ce8FUZ4e3x02RUacY0YO99WJ4DbXfm
zjWgxLYEvCCDnOZdwURiasShR48rYJM4CTNsC0/in5wWuJVqrMfJCEzu/2TkurBb
q/dYdgtcf9G3vkXgbVJasEJVX5FbjoBZ/a/8mjAd1gRyFd/c6VkcZFmZ9NqL7lft
zY2XzcNrEgQhyjdTPXvfr/ppAAngjaP76U9ed4fpFDGBwLA8Kl6Wm7d5Hl4kt2lf
NrmKts5BG6+VxczEpP7BYn3Qecn72j2mbTyBAXXlXXPIAWLZnO6oC1i2hP0rbeTm
VbKPoqPDGfJTRCyqIG80Tr+NciShf6507Myd2Ysf3CtXsQkBmaTzk9g4XKokQNyf
f1HQlGqY9elL8nkQcSesOoSUTf6jztfLkO8oNoED+FH6/NYPMXgQ8MmhyXDywiB1
MQ7wyzsbqJfCiT/Mv7jEGUAwi9mhf3FND87Mg1g+Kg2W0yS1aojDw163V7A/+AGe
5M16e59AdT9bmEhvb6bnCwAY34AVYNviPekKqkhbkSg8dKAdAuaBrUmBxgurjWR7
AXqEoq8d1LN+LN020gpajNskGZMw//HCqUUBpaCih7awl/Ih6KvcpTd9v3XP5MKV
i7n0hQHD3JFTWnbY8JsH8xezadiT2mUJODRfA3YXtbB39bI2pq8CNDx28j2mKdNB
5GbYULrWBxttYQRe9Lr39Vc/ZPIIWGErZBsCv4O5jctLQgm7vb/CrQX7K47tnfjQ
w6VA/X2sTfCBJeqejyhMZb5zSOwsd0UnkN+BNC0Q9BY9s9bUmjovK5brNcz+0OcA
0nbt0Hwa1TrepxowlQ3hvt+XljBSwyuBb+VH7gQQY5q9b//8sovoJlZJ0CG9q8m7
giJVoBQpMMjhvNh1+CB1gXcdqBkU48A3ihqliuITq0HCdVfN9HEG75ditNXsaiPN
GK22sD6p4Q7LTff2dnzNksPvP7oaft115rvs/z2bMjPEHzttpDRie0A/5HM3nvoZ
Gf84BwqKNgLxJ/WO6M/Tya4BM01eT3M2dYP+vuB7/YBXZaRJoqx9IbF1aGUw181i
0TPEFp0eJbwkJsxuIikbz9jMkvsPz6gDp3vKk8P9HwaMvFPLqE2nnEkK0lW7ZSPO
qD8EVaXmj+MORsPlGxjGjf+FuvRZ9mvgMitDjL6y0p3yI1tVupf99A90FMv8XMMm
+sD9G0NKTU7S7/QIQRE1OpxaWbDBuA7HtDOkrtZfWxvXATUvwXa4X9MKzfIvRQOY
l6iuCCFcqVUHvVm+6ZJnj+MVR9dV63ZG7et5glLcQiFhuW1IVAGrUQtdXoZVEOcj
xaFz9VKgabEaJtvXsS0SttKDDaiz+FflKpRZI63Ue0F9eUID5unLukqbTpTSlhuU
1LRLEn874RvJMKTqxJxz71HWxa7ExvJpxII8sDcLSJNS9SsEVYcCq/pP0UNSkBJN
AEkrMDck7jhOJtI+h8QJej3A6kbCnW0np0vQ/k64ISHO3oo/YZkYfSG/k4SJMmVF
MQYPOAoOQdcnQ13D/vI7uuoLK/vtZmMApyZvcQPBKJkCf9+MaoAQESF3pSIBGg0c
Qd6Twg+3sw32lWJpS8vbhwrAJsASguhbqZb++2kCGcnqffx/HrUI4E0G7oI4sXsn
sLvDtVHf8hJle6wYQeAyAxuBK1NoGAEI3Eask0NMpH6bFynwAxX5OKHa5yMvIAXp
2469U8yIC6vjfSyASghEPWBNRKjKfCNqip/xWMJ8QSk4YnR+WQELleCw9Rol8KrW
bsD25puSgbyG3jnhQmzY/ENPkrCNrrhCLMKeiIXclrBLOHelnk/9SfUkj4ETgQfw
4m+OqKuxU2DDKouaNcK7Fagba4PHMeJf4hiEUayx8xTyUJbBpbC6iAGXLjWVx7N6
WapoIwKwjvhaDp09bR4Iqyk5eP+fsBG3X3IespBnnAnww8wEqOZXT4a/6NfAa724
jV5Ckj3V1SYdhuOd0vVvNRHC9OlGGe4jQh7Rt4FdTtmqs4VjfyvoyFUosSFNbZV8
aeXZGniB8dApuABe8Mdvt9rvqJVhlwUFLdaz6HzUf4KrpDU3k2KvY0WPb7BM7a6H
+nfbzcVSb3mB23M+xo/6rh4lc+p8PdnCiMRlGgkq4e/gDEPWYIjH9TLI5yjr2hHE
lMN9URJ36QzoPzBFQflqaitJU8ZWZ1di1p9XsLDuxo6AwIEamBvCxJxS5fOlOIXS
rjJnCo/ex/c6EuIuUnBgWfgFNJsSZ8HiOF7ClG+Y7Eg/TY/lUydrLYFfJV7sa9JH
Ij2EegSTkPsBKKdvRkzPJIT0S3Hdjj0KrIuyWl68+jNJUgHSNih2wh3NDVC0/rst
Iqfj0KWvlFReKrCbvr5IpF0KOrWx3YxBIa3lTRe5kKZzHx3CXUjgoNP8A+F+vOoP
cD4wLL0NWIXkFyVmUyDJ2Yo1b/UY/s8i/NVyb5wauLQpblVqhMKYxGjIucmLRbm+
832xBn/0OrKVJ/Qtx2xe2smidYvUWXPX/eTYAnrjUsmYk2lSqZxwhjerb+q4WWah
CKJ/r8q0ghtiMQDVMrx7dA8IlCzZgFTb5KDOC8MfnwZJhHVz4OejwoqClK1zZZW3
7OJt0CWjP2gsNWGvk6J1o+Srk1VxFXKt5oVYM0GBCsQVmgJNk1lqEiRx9YjvokM9
EoiNRXF7QFCxPx0nLOUUyuCEzQzvnDnM1qiBEGK0dzD4z4MMtHQJmqVTrApZyCfC
JRMdgyYcwagtlrLim1Uh46VwFKraoeRbd2uCPp2WzO3XuaLoShKlKTTd4x8oJ0Q1
yGyiLsDgNMEzRc+WdQHF+4csbIt/Ux7FPx0zgw85HSyid9lkiRp2TyaCDABzDvto
5rEsrB91Lte65VMoSkCMO2GjtXW4sipzzhSfkFIkCl0//MEoZKXYMh59MSYDQkiA
RrOTanIGZmgLv5GVAQP1f3CICOiFj5VH6EHklfZdSmYcaNtpKzVWSNHSp0Zy9FH4
ykgDbn5URRXF4S83gyTrZvnJnyEWFTx5qbYg6cq1KgqUNePlDRYGct8IBGOrrBNu
/ae6nA7iIrjgNt2sCTx8q+pqMjfMI/Pss8yxiMw/c/+7LGavoJjZtKkuWIvqn9eK
Wq7amT/tUl8v6ADTGdA7bEB5CBE3JdQgL6ct3ue2EN50Je4nurKXSezLBQbi19PZ
TFowhrrIAV10wvN6efNVguKbyBY9XwAx0Tgbcf1P2g5kIiUJHWbIx+kVZprH18BW
Xda7UkaEJPYsgCIEF8OM8JNO/5dTMe4BZMKxJw68lQdU0Hj9lmhC/JlkHPgBU9ED
CAGR5IhAqzuIoHv813vkDxiUP73UwnaVSnqxZD7YrZBfIZcCKsx/bQksW4fHM9dy
9KUkZkOudt5eid47gvFQ/yV1J6Ko6thXK0TCuJFYV32HUVG21NBisJQXxtSzseMh
zBV08wPGrvhY7T/qRrWf+L31Sg1J6AMyVXCC9KUl3xvEUYGF9l7OYgTlhCoCRh3J
bPw+J5j3/WnodE9kOOKLoTrCmi4AF5vMji05pVPCZqoByPhp/5IovM37NDkat0dv
/i4A7Qkrn/KN+2AnNsKZpQjeTRIx1rMTtMJharzzzvbNUbSk3IDsGR7KEte7xW9H
wUu0bV1XVy11XL8XBc/76LkLQytvGnrEswI9ryF4LJmlqxvl18whVSooQ1EL9Xh8
CFgp+kIb8VVG4l5luQQ0AK8TSP3d2Af5wXydxIWa8P4nKOHw7lNBgy1qcHBmIadb
Bn4vVAEW+mA4jsFVwx4gagcjMGuZH2cUFd7/u1Rng6QBx+swVUz8/pTY+Kuskwc7
GNvZs6XdcszjLjir02wBiD+F8/V4wm4ww47+CzrpTqb3iV9+NVFvMfLP4Q3yYQLH
yRQ9sMhaz/CizGkV4A1vDmA5pLRtxFYj0bV3PxFql0VROWU2/buDBio5FYk+7G+F
vO2c5LkPAz4i35ibDa9CsocIk0UpvY9eMLhGeosMC1gfF4Dk3tDllcBclDJiJdJZ
3As3KvJVsqI8ubciwm5hUpdIH+wtjFBRxrby9whgufOvCEqEIweiiiIA3QXZqMlW
19B0E+b+mMZSrj0O2MherQlzxGESg8gDEsxeLPnKcGIbaUBriVSbJwui8Ub2StxF
EVi40bbAvxXoWNczPy1lvDIKbaPju6n1b6NNrUCswRZz0VfQAsY0fVkODLxTT6G8
Lu9Ca65GrsjpDbKL+5NZ5dFmIA8Dj+7ZaxjqObPEogbl97yFyOUt/4Ast2UTw3UJ
y0JBjFe144NVDBzRZPnHjvv3J49Kc1WxTESGeZqZQY6Wy4up4B2AQ1ZlONctqSZ4
aMDOZDLY++gOW2jqrDSBQY3OtwtxsbGuI7Na1JGe5fuIu0+QmNOkDq0oL3IFiBjy
zEcXPEUvCAOI999jP1J+DhlBSH3q4773WtKk+EpLnLDCB59KSuKX+Zep4DjLj3d9
b4aJ30Al1nwnwCSMkfNYKHUhKIROwF1YMC04atEt/OWc1bocuTtyS+L7TPrntGQU
5U7V/G9qwUDs93G5LYgc278y9DTchwqnBLb76/WCF9B2tSJFCaKtEAowwiI9yco/
9WWn0tHLdWQcMMBmJuulnN50Yb/R3FRF4caN+s9xzfjpwz8Rni5zHu+s5GyosIbu
URTaag8HhBm3Mo/SoMawh3lns9l0SKmf+ByMhROL8aXJVMwO7uXE7JClnONxKfrd
2WXDG1BI/unAZtwX47cw/c4aj8Vi790cdeoXk706ncrnynbgDbPxPuaSV8LzTw83
hBOmgtiZIg7r/TTYhpZxbJ26ci6pzOr7LSwbekYOX4mYWvPwLtcrv1k86NfmUUi5
NnAt6/DquG9dx2J1tBH0fMGR/lB0gaVg/qE4rpOd+Om4Oy/jgrk1v1I/7OiiS0XE
hBZjRW6akL9ok+Ujt59yiFZ3rp6k5aQgbBInMpfuLOSv5T3z1U0eXPw7Iggl0riv
gO03ldXfJ6TtGKP98Oz+DCBPnJtoFvcZFJsLNoIlzgc/kZP4Tk1tudGu+GxM0Qqa
LMfaUWa5ccc7X0dkbnoEzHspFpEvtHu8WMwtl9w9KKUVv7XViF+YT1w0t88qlGEu
/UCm1vhToEym6WcV2FXG6m6pT0M9zNrGamjhglqGbMJvJ/M96LFA5r5gxFSIbUOO
XlK2GdvS4lsaJ3s8jF+ndM5RUiX0srA9+LlSW0XJrqrqaUuGYq24oJgexQrzz3u6
6xVDhl8pWIWxWjQAURKvUgyveGIknfvJYaJbstET4hEN2aD8vfDtwOKr+Kpf/6K3
U9z5+YEGNl7cJbOKU+Id8Wqmm5jsnYfp+uLEKrURp41ey+nj0hg8af9mQscbIzL6
/OqYMoCMGN2qjZWFiIgRmwgiA2vas7tJBu6GGgOskHbUyKjqBMAoDz2CGhU4cW2u
oPl26pBMeLx3tcMAq0iPiW9zqxTgx0iDZHMrcBmlFKG3QxEMWb+9QKRusYYg95rN
pO+wOnRVg6YNS2odrIK0lcqN4b5Z+l3y1hkVyhSuU7o0hvghCjIq9O0ezRGR5FwF
UA0iip2Rk9xD4iakn7Kk+xUAGTNvebaD7orRr0e3xv/iUPKMovPqgf6wNGPovDcN
+9AuZoDRqrjazc8s0qVTcaE9wvJCr+lhTvm2HObmMd8Boo1GgsbqhY0VBOcw8vPj
71lp3rzrdlyZoF28GVDZsBTrhqJ3r4ret39xtvYdka72csiyx/ku7mTTvrpyhSUG
z+ylLwCYjVYOd7bdJFfedyD34C09pWamG/8aIhp0EZ7MPl2lu/JQouu9mouj0Qny
gUmKR9lb0GUsXiZkZQ3IBTr4hxuSKbvVe7e4rsNyu2HCdYaRPcZgB8wGZ2viENxe
NzomrcCwn7nZa05jsBA3FY9yPUOFxNxs9bdAsZt1n89huB24DIiqGagTyWnPByBv
f4QqFVqqHpAizM0rgl6kEpp3UKhT5rP5eKnJzw3FKcQc9RioDeGaBFsOvkpXpbqZ
x46gI6yo6NR8sRfSbHZI/vNl7WiPI8KrXofPsWTQ6YHu7vMuEQ16Tbtc6jzwY4la
0b/NKHORWk0kKfwIm7uZTtQ8VDktSbl5ReacnC3jjH1QvZ71QpcCObsu1IKWB926
kq7r6VZTSO3teUSxke3prEnNnMiOYBjUOgH1o2IAu0lGEkNNtmmTF3aE9wURtjvF
8N3Sd+3YqcgasNWjuzT44OefO3ZgCc8M7RExxo6SzWdlug2kTAHuZi2D1AFaaZQy
YV3xdhenrKWptLa8LuQZ0tJE84Zav5yt1Iuo59xNrIFgc2BEIDfq6fssYISsoTJO
CaLPX6RjsHxzBudYX1bca9xDGzBA5wurjRegRazmzY6OHVIYAfs7b+RbYIT5Avm+
252POOgGVW8PELeTyyd8oRszps6MM7WCqsT8f1g2N2Q9oxoWQkwBzw4a2RZgGc2D
2WPt1SZKml76GYOkxhdU9McO9dvPJeLH5DwbZ6d+BWUAkN3k2Ehz/F7vMt5ejf0i
cxhyc7ypQXDRTxuPkr0WnlBpdO4qHaXpUtQ96LBDf4H6PSdMuGoC2f7eOg4mY83s
cVyHnJlF/eyv/hmkOKD8XzUwGEePJP+CNNmj/IjbFFiFPAJxwkM6SE8kto7fwqCI
2RItcJscL92bwT0hcxf7bmrjCZEqtGl0xykZ3wGbeBpEJ+WTwilmOWLEqKFqg9xf
TzNNNbfDCePhQ1FAYj7MoyERsmrgvjH/anQJqthH0Es7Slz/pl0GNkbE2PDQbBwq
IH4R9CBWmGGyqQ8nbfTDm11fd4WqfY04I9efOe3yhgSH3vaI3RhuYuS0n1r2yVgs
QGaEaJg8ZxKCK02jkQNflSrtRkHV8/fL1pT7IOhxhOUS7alsmvaiIDdc1t04L1in
uKR6jiXnhUeb8hWv7pt28klf1kSnLZcVIIQp/vGYEpOEVAg6uB+f34W0kcHn2GA+
nddEpz4TtJ03lvofbgzTeVgoElA7VHTzQnKmZtikOXyn5FJI9NYSCcA1atVsZ2vH
2BWXGDbbLJ4+qthRKZWVEXN27OUX8ouLopOJ4uKey7BeidZecVHKBhLTr9InFnAM
LjhkLMiEnYRC+IbU62PxP6QNTm35ZdW6oeMWj7m+n6NM5XP2/vxifYaAxSWEFMq7
8dx0nW9yxJFm0IDk9HxhBnINY9LEAvzFxrcJZ4FL4nCgsttdi+I7/XQcj/tyyar4
1gQ2/94AKgHCVzet/9auVucob7p/ri76MesZ5EtWDqsjkbpiptslM+K9VrQIIz3M
7QxOxdlgmjFROuoX9F8KuXcwT53c1tG4rHB9lbyJT2zlzv9VwToNy+UDhDejM1uu
AmAPxBQC1ZR3z58uJiKTosf7HJ4uff/xUw0w2oAZVGyytH+Yu4Bkiys/nrRtzDMd
euxQzy6n+XbT+rzy17/QXEobvJJMI8vZWmbPyWkqutMmOo4eNKuTeunO9Njarbpy
Pk6i2O4H66ah941o3teqAENNoP4+AFAPt19dsR11MeO72XzYJ5EN/33rBPIAiQcj
c159v+g//X9qaWyRudDsyNO1CyQlPgmy4AHMaNfnqau2MXSh0+LsWX4Hka6Xrb1Z
`pragma protect end_protected
