// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EuTU5Kt6vpGCK1BzLVNPtO5oMe2L0hDDANopLjoHkZuBPD8eKrP90QUIsH6QVHxk
auzXwKSPWjyKxi00B/wFYvP0XFYlp2ACBdUeJbLD+vObWICl1D1ORIB+Z/qjdeN9
Q9pjgAKlyPw6OOYcJh5hIb77qiTcJEmgg8x7uqnXTao=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57024)
ia5u55n6FkQEzWy+E3GCHrfnczWsa6r4oJfzV3BYK6dazDVkG2CzFsjdJvjm4j71
38tSfART7ZoxEs8omHFHnJM8a+xrAF/PDBOQ4k5ITQW4GJZn76S463G/mvwjiL57
uSrCQA7ng4WITVeq0x4q6cw2cOxn+pOFGDYNvktGIgw6cE0pQ7lWpzofjixeaUXI
wtz70MIjs9hYnYMLTzzY/5op/wp08dHw2GdrLxm5HPGEhJa4dFG/XDcSafC6nGSr
XaOou3DesLS6Ghhq8EQhBeUtPPvJUjlFLC+U9/hZMuz4819oAjeOeosgMI8vFnpU
vryLaec39ZSIVc/6TENNRLUA2yP5RAYU+FMe5gVgYmMNc1n1q1ca30kHq+KRoxre
HLJRtfK1nkJrLm7wXr+AZJg/LEjXUQtPWpRtR4dKhSAtGUvFVf7MAOH/uRNnLbBV
+4LzdP9h8DZbD0DPTk5W+6uQDjsHF2CRWklxD7weBZyH4eLGQELIc4xkp/0M8A2h
0rvY0S41t6EOwzlyZLM/4pFV8HtUuxkgEH+dO3Zy/Rd9Zb2853zmdX+zfWeUKSra
sN7kf0MAxKMydNoVkhP6l5XglGg/1Yv4/K4Ybcim8hETjpYnhmFL3Huguaiav846
7Y+muNUBbcandMGb1jhjVY2FNpqbU2fzMMEQLY+SsYc3n2x2ZBV6lOy2MCXS+cfr
YDZn0/twxWolfzdDPp4lUucV7ofnVKtpsqwrbVwQwAF0VEgNkUf6vXMMlcgTm/3h
FyXaBogiBz2M/+dtkZwH2qWVqk6v+zth0Kn6Mg25fOst8CDBCG41z/Uomw1Qd7OZ
D2s1deLF5w7bRvkutCQeUBEaw5jyZ2MXDCRyVj6cW36xqCvtndLIDeKsSMvWecuy
SNVSefJFNU+fQ9iDjHTuLBrneXt+Wdn0xTaEXNCZ96VTlwho7ud+vvJiVzD0NDKC
R0GMo3xSO6u6jGQhtoXubdaqWWf6prvbJnsORYlJZO3T9UHb6/4Egwuiz16QKiKR
3jI25l1b/uzBUJMrU8vA3uad6JsdgQ6hrfP0LaRNib7HFbEzVIL2r7rtjsZmXN6i
3vTMa1PCTTm88q7UxkBCvwCh7MJ408EKKNriHOxLPaNUw5D3yrDgUpiGvB4ONbF9
8/Zkzj7WLjjydVTMV5KKY4KrFaXbgC03Yvysjmjz43NWE4fdl8V/ZYjQWALqWXMP
X+N61HsMtAM4j8iO+kZ5mOLMxAn2tsPN/uhbqg/pGGbV3FWTwhh81MigeotLNEEV
nr0MekDEffK12AqrEMXwYlnCXlGpIxOLzzadysPqWJ/jbDZh3NdVNdQBYDFJ2jki
dJpkHYknPJ9vvAyzT8blMYzQvmWKJXhrdzKsZCu1Rpvr40Gt6YmdF4eUHNb5DpvH
heHy7/iv3+GuGFKGzLHCGYzwz4tqlena1Z5Ur9yvKdMHKdC5HpBKijpD6/2XTJKy
C820N1CmZnvQdxb321ul3LGqX85B0JQZpngkYUS4EKQFv0wXfJXmgaJ86ZLwNgAi
3CR/k0kThKf53KZJalKSK168CdFpx2ci1rnbLGY1Ow+6NqkLeaoCRGmqRtFPIQiG
wNs/tWWJHXMljV97OODYu5DInQy0EicCpuo10l71zLWnkmFgMW6kg0QMC+RiNdkw
lCqrG1F+PiYQuKny389RVTHIeTW4PYlT2MwQXv30f5iZZULWdd7BglQJMk1I6l6F
eGsEtcxWHiBVocWQFi7KOrv5AJtVk4NN8j6efcd4PzKUDxXfh4+SJtGrTy1vjPCD
XSaJldaDuvTvJiconulSBxbfgtBs/n+aUlVG++gcytg+2LgvS5LBObFg2hgdgJaM
NN0OcYeTyTO8TU169j3QsYgI65NNgGq7MLN4jEB+ojkYn5rVarAsdkpvyq0mEmpm
4iorYteBS+mqS+Mm3z1JayeYDpTbEID7zLWOU9UYxdZ0fHEotKnHCjQ3Mhdcsyug
cJ6JrBmtKdzwMSX71wAfJyZcOpNBDlJR0pgpQ3hufYMW0HKWwPu6ObcbWd7js+/T
sirHDfaoRSquOTnpEYSOkttIm/SZW1azDlffS/vQlrsci1yNvHOxpj3+ME3jE/Pb
VRoNmP6xA0RFpqHH2MQ0ueKovO2J5Jam0AB+U48VPqxsz34r9aYUQNRL2eW5iCwC
9xheZOkenvbhhs1qtiugplFbZrdcxPaphB5CMbadq+ljgPldsnlVqlNl8aUMtY+b
8ioUXVNXQU/WPuhcwa0OB8JCDunzQi1HQxGk4e0N/hbHuIfGjoJ32iCbRjewu6dx
cKWBTVg9uLa/c86aHYC965M9HqyTBZ0ellpqVBl/hC/wXqhqoTaPDrTThi4uCBFA
0WBsTy6MNtNjN/cSbqjVc+bq9pP2UijFelUSlnuATfC8zJ8z0vPSFf8FLROQJUic
bbxbLE19Buw7WukVQf2UAl6IOzBweFX5Kfww/KCTDjsT8FjkrffXgp11zdK5Om02
6tlpCb9GMxozvc5WBTYH6IclPHpb4QA19XjSfyNQfYWyjqwcjEIvgmwjKZM+JdlI
ly66B8+I22TiyHe+SS9zcGowpiP7yM5Ovcr4LFuBqy8ukgRsqa9fw4vpZQHv45SD
1nMVHgTnh77eWCkYXf1gh/52pOqDMWYsFU1jIabGAi6ElakljmavLi0WK1VjPpZu
YesukWIa7MaTPcpbn81xQ0W9TjBbmp2EK/jRLqdnNsXk8gfiMTMWF5fvIQR2nq9w
XzBGAgMBbXle45cJIknUEsxl4Yi4KwsC6GU3MtKCOsNDTluoaoh4umkmuAyIOso0
24lLlM77o/GoUwi2A1FIN+dCTw7Uc3rqV7OV+5BevvrD4j9W4o1dUf0sQ68PmJeN
Xj+OHi5rRDU+sY1d00eXZXL+mX+dJynHV6AS/fBR66acShYVzWkpVLc4mn/xGnWM
tsTajPIwyS9dxwwbaC787ugw9vI1pyWefCd/bxaEthSzLFWGQkpRPmoFJhqXBlCd
g3ivu1/dkEPSzjcUYL2Ay1VzZjFYObFkGKQ4Uyly9puLMZFT51qDrUuS51l9H9CX
Qdc1S+v5/Vz5rRcISURMJsb6xnC33MCJyE39gGnxJFoelpprTeJWTleTTtzVOtI8
VwJNwCWQD9d419aX1UxEXRRx1gPMmOHKLs/+enWR7VA5xwwfTFGuLvfP5iF5sLgH
UtYSrtkXUdOgUM/PDDb2ADavJwvEgewcHHfBB4lvr6grtD1865oySsQRHoPFtClf
4lct21mWn/sdUdgC2x5MqXJXCJ9lJQz0VvjxKe74prSe1vaSlikv/TUu+S29lzrE
wXWrVwIcCmuV7EFKXjFSkflTwjcBRdlTZ64Yzx47JQjFp9bf/BHrPKhzLjAzHPVv
VKdLOIxia0KxClKGzUdLZurrM1rMWW2/yrhqYoGlpIQT7fo2eIjTo1JzR7s66Qmv
feXHUD3GzVsGcBsYVvhXLg8Uw+wYU2oxGFalfA/Mfwh5H7dCi2O4/DDS0tuVOgT2
Rc7cLJS7syzaeiLvyol1WAYxnG2ZQ2O0kSM5t10tiXnsBiRh8ggdf1899zBsDa9r
mYKqL6LjHhV3RuRPHS+7Ah5qNxA6B4ijK0bHf0MPVz/FIhZWmKgjicn8eKxgPk0x
oJ/qz0UC0isliq+VIrV6ioO+4H3T+psLualGztMGnEGqEeFeUcnxC1mWdm0gdS/7
yTowerHzcYcP31QXkA0iCaP8RXeXzJmZTHjWtVm+HTZ8qK7iln31HrqeCbjVFDiX
kD84pItagzN09qL6pNxil19Bn1fZM25yIu/DEh7VYiYcIqSDpONJC4N4Cx1k7wiE
Hb8NQwyeWGDE+88mrB/qYJxdRHYWYxPbMbmc2SGZh4mb7p2D3YaOcdlU+h4HlSzL
uMehbBZ0n8YlnvLtjEyWtRnskmcsSxdlSohG66GjeejjpKMC4RS0PA8FRgm3W/eE
FvCU2MZM2OoHG06wCP7XLqiQS8QJ39tUiMzpn7rIPjbHjncIY+3mGateRyEpQVDj
NMvsYZl5tGaM8/Aqpx/Vlm7qDhP7CamtaTu5J491qAXjn/VGvh4dOy/DMikTpVaH
tmWoS3Pe+5ZOxrcf+oZv2t8LvreG6NDfNkJPGZGFg4+Jel7yLDzYR8WwyjMBd8EJ
BQlwr/Uh96mUuHOXxukm28j1r1E03dOSQSirRZTS+MCd7txjcAi7DcXGCuS+oeN+
LF+8MYL9Ta/b4Ck11Vp/jwy/ebsrQOodUdEcRYbWIIAewLJ8hFZAP1C99YBbx5+7
AOQ0qhaVKUy0FTRyeXZIZB+OgUWQLIv61bINVzcHpR+C+o0w71OCkVKugwwxeD9O
d28O5qilzk6CmquJDvy+KtJ+tuN4cUKwycD6+fiLwTkH0DGYC3DM3R70Z9S0WQvQ
5f8rDWgoV+J+iMWpwdLGRuqpN+vWkNH19A18QmISdjSwwa8fZZDeog1jEs9GCdpV
MZXiHKJhVyNKrrVxvI59NCO1cyc28A8pAvP2hHKE5a6mHr3G8hdTrUTz2vxxjClE
2uVecYM1fnHShr98+gGbAzaGbU6rgq4KBTAj2L5oW/HB032kSyL2/qrN4sb01NHX
9ZuLFVoD108ZVXWEIfrajITqcfFsXukoTCzsyipsTrR7W1KvvN7XKoORDe+wS09w
E+1Ao6NhbG4ZB6C6WGi0yP8bR+nqF1IDfCZzunijUMP3U0KeRSGMWojd3W1uedyU
wZvAgoEOWChdo8PGG42OL8Bs2PoZv5i3KTwJWeMLMmre24qslBsENOjIDYVXMw2l
U+HuNmx/XgUDsyjNGUbrnSyZniJ7TvOWWyzTJPvY/2t/fAa2HhprMD1c0s+g4eCE
WDKH0qAWFdRDBr6DJ1e9LVba4cSYeLW6Pl56fjMoyhd/AHs6HJppgOX6nmw9X7Lg
jPfkcPTu9WDm0T+tmmspeRqRjEIrSgqSkeI2a5XRSfs7AsimIdy+mEKszU5+4mro
CltIRtVbmvSfojnFzS3XxYFeOdEqYhxfJVwjqRWVmvFis59n5Tg+Lu5Aza8n07mU
verBSao7VvxSK4onDOwiMmFuzm4ZRoliyfy7G+V0lFYERSXTkAliNFUOpO02dfB6
6o8XhWKF+Ly5ZwT/49Bn/0dTYR3ZwziDbDaJ5S7QZ4nF6oYx35JSDuKO7df1R7Kd
XO0qmruoucVkDnTXiEnHDWIcwSJw88Bi0iCG1zAb5RV5MwVA4ghhIneqzlIRNjvo
qTBqTxmfISgGrXI9VA3OI5nO3j/RrUfYIuzsP88cxMxkfFWPqrZFs8y3PFaNL7SR
63bUjOfF/vIbTaHnlx40gZzgSDWfYXGlt/f1Dom/KWVL8UoBJwGrgWR9z6NLHaTf
0umlczILTwVMge+cnNyxOZpGR3jebycxV5RyTgowc8WFe5wMAIhU3CfMky7kobKa
x2QaUUHM7kgH38OW03uGFJJT2M5Asf3LEpVbZFzfo06KesaBnR9JEeYkZndS1Pb2
ipEzmA9b7pw4X3x/OmQMrYxBNgu7S7JM6q0UnsTkjjcjL5a/bvHr8KyNmvzEyqtc
Ri5bS89OxURnATcdnw260BnpENb+BWyEEI3KqSq5KnBWn2G2PoNYzMnJGgVLon5s
UM4ZMVAATaioMy7XhvmzI4TaQ5Y3dc4RGT5Zfvn2okh1Vc6GVqqDL89UH/gdVlDv
7dl1HRhplCFZrFJQrjq41A/m13cobmJS3SrH+cMFVy0dqtSTHtWCoqkAJk2FVl8M
QXKuWxYWiPNHLbRE949wblLizQTyNvaLVWi3EYoO5YkTxF4/oX3keP6rxeCLhbm6
WxQTXTPZxVv/dQH4flV5Qajr/rxuWJjkVsiIp5ls3lmBRVKWa9wrTCOouIvVtsjz
yw2DhGO1ldrw4sh7hNfthmUCd6IHy91vLh8MrDWrD4Ps3ONqzvye8srhW+Z1C3pc
en75+q5RbOvA8Gy7Fy0X0p45kJITQc+VSvcf5jn1jhK06Qty8fcrn1aRWHFtjZwS
/q+NejNefXUI38GrDfpXUtrjRg8gUu0o9YiRF7GtHDP+m+EbxrC2BUywvH6Dji5Q
7J2ErC9ccsWJpuW9ynQ/RYEBjuGvmGjUYinfhX3xf9Cb9laXBXMGuPVLjj+cZ4fv
tkmR+IUu2gD0jluBIztilv7G9F73OKzjYrKosCfwnMjtSdmHDRcrBnO/SswOAXjm
ZYfVlVej4Gj4lGN51dH1m5FVB1Iq44Z6HNw3kN4Dti0qo35Igkm6vSR96gMzJT6H
AdolD9UajDSn/B/HEAS1LhN/XS/IdeaL7LWYbK3dofCqX4JRH8hoQ4cylFbXidH0
RiAw+9xKhbCegYr18Bg9PUWQO8zvcQUNxIaXIqBn3nKv5qZS4D7qFX9Jq+G5I9yy
uGAUvWz1K+mpcFQK4YSiPFAL6HPMS8PdPF54wXCfokh0QaX1yrkAPLNCcW9oDt7j
IedjSHHhXEFogyN/q+y8R81BaWpgB0H446X5ORN+KgiUa8++XpfzYHm/td3nfiMY
ytFTw+1xpy06i10Ho5r8RTmcSfzLiHydVfQBZcS0xfOJsVDtre4xvuOFUlALYbUN
W6rFLtwy6BtPIeyD7PKoR9p+rS+JOJHG0FEFnQNkJ8D9xaHQad34GM4S6r2JIQaS
t8x8sDa7A4J2WW/52yjvsFNt8ZbgrduQOmjKbsfxGrAunwW5JW3RZYcaNKnTASCb
cAzXUM3LvxPl/gvXSc88ONA3bFzg9XqwAD3/1Y/B0yzTWLXLRho0vPL+J7W72L6b
yTbBEc9vq98nVCxsOc8LcfHNGKJ6sf8DFaBRwyLeBrydLD3n0bLYdCQhWsG/vFOR
Wsu3G5OmRQ9OCbQ6q9WIza11JwbwMqlRFQIhQGohSWe3QEBA11WgL5i234N27D/Y
LzS7sWpPUJmfxdjQyunDjIqm/VMlNNLci87e5XaSk0oopCn+jrcLINdqhWQD1s3A
oNH60/OvrNd+6gopNzWpljZsZDvESMBKEtvut7gVvjAc7WfiQKsbGvU4jsv2MoxR
11b8ISuCxMX1qEfRU1gvvvI+c9pkIWZ5lPaxi+w8vCmg0jZNoy6Y5O5kW9/r0FCF
FBfvkdVFiPv8j4UBnZ+6JFom99j1TWGgK1jFJbPDkAvYbfD7gaP2WrF2gG2ZaXSL
ZtYLPMeWIGckhNtz4NQ0UlL+cyw856FtEUerj+bTbYHY6uMUMiYyw9752NDtXNGq
Bc98++TEAqr/5TU1z4nR6GGgtex+obBdxdocvGYpg11nOLLaxdhT1/mCupxGVdc1
gfgD5S4EWT0rNew8cBH5ypjdRfydo32PAyOEFpqeX7NMZIAPAwRjXYse4fulTuGo
c7ogJkXI5Y5TrjY2/NYn16CJw3MS4cde8hEBQ7+wCCHTmyseoP4V5RB7AmwOtjRd
UJmplcXdDIaKANkTgo8oU3YPx8IksdmGfqK5cLlUuXGoZDA1MPCXbqLXDTKHDcl/
T4krix3efJRdBjBMA0unDEge1lW24FtQnaCwhP6qOBx/KILPqoKoG+cEqiMLdsbO
SF1zR6CdfBCZKt+o6XpMUVd1FFHGeMOol/zEtcW7nOeCEGTB1HVEOgil937iPjWg
vz9/MR9g5dAC+Cc+CNHgIoHWZ+BsopnXur/5E5qGb04R97caagczLkSdZGciQ+f1
yvYEr5qPtYW49h+OX7K762CZQgARBWuiIMWni1H2ds+nVnRBgLMcjugAych+HkNM
7K9tMqTkqRDwpMCxeGZ+oly98LP+Jbp/aUR80CYdyONdFY0fXlx2epTx5SdwMTs4
QC8UuWBnLjXBnh3AC06A+czADFCXOm5qQpe05BOrY80DRRuMNthQ1CJIRlseb+fN
hiATtk4WYTRImZy53MMtpD0VokV25AAAwAjyw9SNLkb6QkXyGTxpqLxllWJkeIOC
eZdnlvFzYyyShrfW+R5CcnetDFTWUPYvE/9XOhvVKQT0snKY/cUHe//5T+F3EESH
QWpy+HjWxkchezmhnpqFl47sDkEpHUojDvVXkU0nvH7MZpZFpcfmn+uBE+ndnGMv
niaQEO8dJ1uQeFXjlyG+HbPdieQR7QdAnonXPHVrvCcG1WZcdDgm43nJI/VIN6qJ
fXUQriYT3GhhkkjVEwAsHZiT6ZCmQ2eOIIS8pmKgNnlJegYyDRBB8AfneAiiPkr2
9elKm/9ybDSYJoxvi7of9e8tPdoXnxvV9MP3BADaMCYUPygPe1Yjze8hKYtapgJK
mLxdz0wgrmFVOUuiBV4kgjkHEcAZIt0QLq47dZ3kTTkAf1sSNjnxnbMy7yAnHxhh
7EfGdfB7usIfrGN1RZaWs70dcO5XRJRw4NMn8UNUwAqzH+9knXqnrJmAU35+UyJB
eMKmsa7zXHwoE4HemlTTEC62pimC6tbQYCq3+7VylqlpvkztYYZnTYWmtFUCQ5E+
KUuna/9TeLzkwACi0bwUS2Q5DL9Qvl7d/JpsD6A/T2GBak0GJr5c5x+y6M/nzyk4
SNuAvoQy2IstYJS4TqPUxP0nuuzd7VdcumZvnyv38KlSud31XH8++CxVIZmsQ4JM
IqRwl+F4ZHmhLeYxdii9UN1nE2syQH8+I9lYCdfKjE0kqYjiYDTJHYTkEhKLVAQg
7XPw+5k3Pg7eezB7Eg8x4hhUI1EcWZOAammyO7Di9VBtOv836zSrb5gMd0JTNdTf
56ULGoYJooyPDS6cRRzHcps+yt7ax/7XtcHWsZxn8kW6eZcHSSeM7OiXpeCbpM1S
Tl3Dw4cKHN+NDEaDTCJpj+a6gann0cRHzST3FXEIFVFV/XrxcKDwwDFRdR9OkzFB
3lo81bA0zoli0r1LQai9hvWU+SryS538G1ZhIKu/IT7aPM1TjsGZNEsltnAqYcgk
8ILQn4buEX2yUtsWSKcoQkQ4Yw+cL0nzsGWoxB32FjSjtHm/x4OPsQWs0QY7+yLS
9dVD5396m9AEpXorSX1nZHArDTNIV3Gb8h582kKiPhOMjFZJpJIz3cSjnAFq9H9L
sLxlmGuPx01I59ZwW91k185VUXuPZVp5+Yfhx978zyUUykhpUOYidfh9qfP3NDeW
yTiQJocyxzqWSfUqNd7EZcvUelh53ICPEX0IFMchmU92hxsehh2M43Ld6uO6zhuE
2/k/oul8ogNdlLNNOqQvxpq/Hl5KOU79FmRgpCORNM1Y80p067HacCEpPKPUMSjF
nsLnnwgp6ZRnQFlksbDrlBwqsH/Xvq+JxzdKtavQ7J8VnL5GZCBmEdSc/kBb6jkx
1jle7Y/A7uQmx3t27wonGD/R5/yEWC/JF2zMwBaapFJZTrNYwOgbtWZhr8h15tUm
PV7e3xXBrySO/s1lGTjfSL0MtxFLes9/siAOSyoYfqdlgPRGRK91P6aggrTiyFIs
13RLuatQvv+fOznxZpFsA/HIDHnSSwgPp6ftDdwanlpzt5QvCtzmZUwh9UpolnAG
WHgdtU0JWK+yZmrI4bpMKDlEJyfUsriVwLMUReGvZT89IGKH1PsavFsVeAEtVauU
QiwSYQeRBy2wmyjyjU9rdmZnii63LyH07FMk9cJtCFI3BGNxNoRvISkG54bd+k6b
DbIJ41XWxs2udklLLciXKKcokGr9D8bO3xab2EzOWmNi1xnsLuWPQTe4L24ApgQF
kYIFi5hszBtqBzzhRHLmO8zD712wCAgR1Q3adkV9YG6RovXMluqn97QUFypVJITK
8cYlrnPjCxLz6vL0PGuDKrv2GWd49EafHPbM2MCHhYXVop2GI6CGMEMpjepuKIaU
+EKw8bMrCGC9V4sead1hNzyblue9RQ2CAaxeoF/HrXTi/LwC5GI7hm4Sy/MwlPT+
P6MA75w3U6d3y2RWvPdoqrsluDLXtpKGRfQJzljVat/mrM06my51rOJpGEPzF3X9
rqtAB5iogPKMPxHiXC79TO8he+Qprt9pB0ARDNQWeAFhy8M0X6RcojgO+s+HmTDw
N/wRZxm2gshckB/9ujWKsrbapaX1C4tcWJUFirWJa/LbavQr++7WQmsJowsws/wP
Spj6QFg/AdnFBh8tdiPUhIKcS1g2KLHsvabXO9VPxHLuyps4RkyWuQSs0S4TNthE
vPGTRFwKXFs8X5I3tg3Z+lf144r38QCV10W4zFItaGpQJ6bHojwzbwCLZX8BIJJG
fpWmEMtDXq228ReW5KGPJbZgdmYDnKFBAQq5WbJfz3zdMbqRGCUtyAGkoePpTQaj
Oi/7OZjeFDCDXlzjeDNIW1gKICDBFGLZlkN0A7p7GAX8oz6DoN8B+HYKhEL4PfYA
QSQrS1OYi6qmhE3Dyq3q25Qr3SsR6YNVpcHY2MTXmMK2Aw1x3MzcVRVUPCcuL69K
MKyGYaAqTjaBu35as4W0VN4U7GWrz8uzDhrxHinDtv+gSuE32B+vh12X4k64D8Xw
WVm8gZAIdm1SYM7jat2hYp2F61lmx/SitQ3zggFz1OKZJ+TLBdoOCjGDWWtNg/zh
XuBlS+qvIhxyxwuMQrBaOK/EnWXHgRJ7xomUmlQub/vhVTLxPaa+VhNYX+nR+Q0l
Ub5R+lIdazxo3gq38h/hTDwp4TWFrbJgpmbBB0DLvQewLTYaF/YDYePeKPFcu6AB
jpzXLA9gUk1pM8ypPpbz+DeknBI2q+ip7Tm/XUr8korHpp6Q/vkP8yXauWH7/Bhd
Sn1+K3p6y6aJnNGTpKOX2hnxmuJ0H8WPJMpjyZPu1HlQl84Gn8FxeXGHfJEQqJeP
3d6qb05fUr+z/9Qo3AKV4O0S6MRQmAPGaD5zTa/Ykh9MKOSq5IeCy3D97QgPf/pQ
mO+qrnx/7egqtyP1hrUW0EwvvZOxSDIyxFPesvdxDHspacvfBw8ayM0zZmGxttmk
j9GzNukhYvQm1+sg6bv1vkjNg1eZSgXrDA3Sr4c+CX/4ZhkeJdou96q8g6zeToBW
ozQYoTttuRBaLmE/ejmLaLWnxyYTMtCZpy7DvNAxZYq70mVy9FweT8hg8kltTDG6
377lEQnqGrPlEEZT4GCDDxdH2p4+RYlKbcPYxXLDJEuiDBYPVcUjtir+97cCJAKO
XnqR+xU9E63vidQt+ahAwvuWFnvUMZikS3b2cCFFZ4rYYgo7fs4fJVG9kqRGW/wb
IxWuvpD7k1EvQysj/0eWHKTxV+wa3e4A/ekl9KBs7Gz2WmVWcy2OTylgI+HDm0A8
UeI/WEjNrCMV/5f8+IWr8tCU2r8UEorLwRELy6UuEY+QrPUtBLgXKyW9T1BjgTw9
7YPTZl229qzEfnHAoI9QKliK2/7FAQaYaWZr+Dr4hzs9PCXIHIFSVXXCeyho+iTC
yqPRHOOl3vVMqj+5uZTAqcZjVEgKKdxS1PQ2cvJtjays1Ah/QFklXoHPXaey68nZ
luR4xxDziUSlh5Pz8mqE8h1RIxUILYyz8FesuNYx2k03CWkGBs4BdDBkuDB/8MU4
m0n0yrSqpnOPFdN+Ys0VAUKbMxynTdYlqeClxLQM73fYy2Qt93LbYMHKS3IRMpbU
3IZqbR6rpJ3QZcWfE0/pbY2KSTnfmobma1vLUeGRBWT6hDyg/Mj1YKZFONAopKBg
/E7iOhIJVZBAAm3lnbFbgUKKCjekG3r+J3f1G8LDtEsLYeJ7OcJXUpxl6YRSHvDv
uOLx67/+5R1c9uk7s/Y1jPCgCyGF2SbdcCXOcATCnjGYxucJRDmcg6gQ9lN9bXri
7mz/w9jvvzIHppRWJzeimVq4Y5FW+RVfBPFhfxUgxmWCDmEt5Na9j+ZsbRCGSK4k
GlpZ8oCIFqUqrA5jk4l+Qof1zHKd8A57z5gEA2C8gD1oxZc/BQ+nUxu7Wwz+jmbW
XSRjo9AJvN/SKzaSRDEXeh/sP8EO6t0u+vQmZgusu/wjwpdwTQdFApqncjy5/9kl
487V8v5wUl9B7j+T0xDPFe+F8OlAA0umvm+3VUbCkJUwKUEC8gipb4nlf3F17ykD
2NnU7d7GRAzldgBe8VJEPJ/SNgujdW1+FaGokcvWZfNYOGWWuHRnFMUPHJdPgrar
xGzqscNbz+gU7Kr3fdsU5P2HucIwoD4tgBPNByusTvRu2oYMsobcyGSQXUHN8prW
yYl/HSsP79khHwlwV+Sdya0mK7WtkaBm3SPSptUKKtsaSrt8zO6fmGt79v8Iw7Ju
Whai1IcjhJdK6JPbSBRcF4A+GBmpA1DbAtHm9HO6lFw8yW26B5XdsR7wT+weFH45
eGcy+vx+JdBbR2sXoesqQzYo4EwXAo8Wyu/ujTdy4i4WDRnwBAtSbH8U1MDA7vTi
UEnbS4CT4IblI/3LFSRTkmgRlhHD0vyh84pPnpzAWLtgyHa+ayNFpZPjg9+TJam/
SqcsLrGOF1iq7qq5i0jZmJEXxfSX2+06BmZ7quizG8b4Hky31zGljWXRf+JWDeZN
gQUyifRAahXy67SppmD5dJd7AcpoP6ljs8ggkceIH+XlwskgTsuSqte45GlgHirm
T5WFnVRP20qppMI7VLG8B5ovPkpYdv8A3yZUc/vTl5KFIofjWc7VIr/W5ELx8AtY
tJJuozWAecF1GtpL8u+9vWPo9J23NzCzqsYwgQ4giDshpcwYZkwT+FJdicRMGIjO
jdJqKcOmtaJKc2m0afsSQzIQryGC/hPi3IdfRd/XbzP8YASaKSVSAOI/Qu0XzIJW
hYMM9jMNazFrv8cOesMTZRFVArJbb7W3FGraxGV6FOZrzYO0Y+KGl0vS7IVe3MqV
P4mh3XHQhAoSNMeTWJLD7HH0gp6Q4FiT6GylwImy8vWjItcXAH3cNOZumK5ksCVp
ep3HZoJzuNe68lku2G36oEvZS9StQNTJNAjdtaG3s6XF9bv6GXr5r5DjIQbCckO8
dIG/NaXsBawPsAyF81y+D4uFXEQ8MSzKgsgtRm0yEwbRYryPUZxHSYbjnmGhEnZU
E3A073Nbe606cELspE1cJg+nIp6A1+8PQCX6feVng9vLJQp7H5e4q9qopssfj9lq
lrHEUlD+CMxpN3JqVuC6CUkzcWY+AAtrM2qtZ8Hh5r7IdO8SgySi57bw89GwZIrY
wmLYybgNK/iHGJtpJ4EhJgPHAeQx2DSugBkwU7S5Yt0b4Dns6PPRFFROdZIf4qyQ
6deFKib/15TLQjrjvM3kjUGRCz4YloCvskr8s74YIIKtzIimHbLUEnBKeuD26zbI
a4xurwOgyAjFxzyykJWOsR6cLrh9wgnjaNb5XVMzk5lb41P7vRUgtSDkHCZpPbM2
PEVVM2+4YbRObdFLCWo3HwCTHOmFYyrNfbkTY0BbEwPDCl6MHsvI6Zg767Xf0gmP
B1vw87apYu1YklHfmRgcIzjig4W695unTwU/E9GLopeiW3+pUC0HpPKvVeHusBnu
o1TrK9oAMnGs+DaR00KWOqCobbyhVnxsrY4pIyCLVJ9uIH9ykAaVvccDXYzNRjEG
DBjm4D9jw8WxMxIATzYMLLnHFKz0XNvb9lDYjI+lMP1RadaeitgNqBh3kRul7EN2
tJUEaf0K94R1BY3oDImEMf2SUsGEmbue8abwsYc0xToBJH1s8DFxELNBxt0NfOcY
cJkLhYmHkrVjZFbsPXDFWLgvyQcAiDrc9frqsaYDHV/6XwlL8b2EGJEVZOv3Ps81
+4ScufT8p3sm8mJEnWmfAAouRbq+z9Tx634XhJ1o8By36fnb44gYuLyEuPXByRgU
Ml7ybtpbJta0YFYLGLqhj99/4wxXk/7yvQ5kXG1a8IvkTX2Jcuc04AXafpnqxTD0
fini+H1Axu5JOxTgYRLR/4+NdoAG+ATjnPjGh7tlIYDRR4KZqE4SOWdN6KB0ZbbL
W7R64sQ69FbTgw3AHfSnaqA6W4JZP4z/afxKX1QtmtGgfFMVppgcuhIKExY5p6C/
BndHox3V/WHFGeiYfnk/pel2OoboNWB4TzLAm+6wsfoSqGXPZ/Y3X/DeE1gsWicu
0ZISpGXdJAjKyxbx6pu2TCUhoKnKXefY962YqD79eUA5qLua3tXCDhPKLvcRvF/S
zAKNNvy5jFjnwWK42aYzEPJdnWLBCyyhriwhjH9zy1rJQfRcIVkOdLYLhvsyd+ve
AW3znD7oVImfoXjE+b4YInLsLMACYPQmWCx8BtNWVQALFPuMdVEQ87ZHeK3c6WI/
dayRGHpU7AfZcn/OCDOgAeSWO22lBhThO5aF8N692k0R65DHmumo0x0USMNna039
ywdbzmackqWsF3dCZRtNcso+6BtDO0ciAITs+H7Yciqa/lG1JpID4qL9xgGNUMtX
DSDSY37uE8HsPGth0pv+xYc1m3b2l/gPRr9q0xwv/2bqwosRVUyPZWUx79GypT3V
s9tz1xeu/TZntNUYMzr1l2XbQe/g17L9gYWfndDAIGxj3uMY0LLNJ+8BGvWmagAY
+Yd5UHWC/4SoVyQWjpTgVofYRNhfTmBliur6ooIaKxUnlXoLHczy7ijiQMtNVCaY
r9b8U30rQCPx1Vu9h0hqE2QaZ1cvAQquSDQwPzHHTdhFeaV644kBFaeaZU3U4YFV
OSf642w/a6Z1H22hh+0AEzUjxHhDk+kpbP/ln6i0KKcS4q8fXsJsQC2vvr80wztR
TyJfanU57CJOk86bLWqLJ0rHO5IBzF5N4RVThUNLb/34Qs3xZcJX1aAuFFVNb/bk
07EBlioOw4ELiQQQlVxsMZTPieTTSFgskc4jayNDf+teBNUy6z/0cOCMIJqgPJqQ
tK4+pGCDvvoXdWluVua2m4SueRW8bCtIqtwz4C1J9Yg0SggQpFuUiobAQbrPGqLq
YMSXqzzU3Mdb/bek5ohLxVV7zQUPKvIA56hTTy6MsdYRGohcj01bNisIuWpy/6jP
FxDaMjBk34tDCwiV0RNrpscrPrBGu/qsfus6RsU8yweNjeYD2/XPKwVPQsu+cIzC
WaNEqjr03Y5nRm9JRSkqW752p7gBEsWmNeZh6D025J8Thn+2FV0GVSFCRtI/I+Uu
taEnWZzbGowGPy/v99oZvDBgs5+mXLx8da5d9mEZFz9UxgxgjwdZFRabN9wvIHUd
UE2GiYHy4bh8dXhDvtVCRktrPXv8XsIeViOk7VvVX4VRp3WkneHIcG9ZV7n51XLo
ZupohLhIX4MA8gvyOGxW6JqODLQ4F6CntmmshuaEq+oDB6m0j02z9JTlkx3AI3Gh
/IYBLqML5qjF5RTA14KEWqANfhJsHxY7z55CtSzcSHAXOmqYEYzosGkzuRE9hWqt
/5xzqU9PiHeujlXNcnXlIdQ+GNaH2gGVNsgrjd3z1jk7e8wYtdmNLeXn1oeLATuJ
h9BXXaPX407oqY+JZ8rhCo6+i2e5b7qyaeyJWFFeRPaD7rCxU4sNSMfdhYXqEMb7
EXh2AWLwbharvsDm+imgvWmmBHaubl3Nwa/6JrLsbJAzBx4bwbkoQNK2KPX3SBrv
bwCeGITNRDmG2DxMqWvUWli26qVE++euAxDYwsNO5dfSytkVXixwOa7kBrGcj81V
ij89of20UXn6HeXUFHASHov2843lbiK7EcrEpLn4pwPcP+hvjam3pQky+X1V6JdQ
g/JtmNa2nsuVi9Ot93SjdxcQcgUz+3PlKjquGpaM7ereAXQZkmYaDv42nH2RUjHy
YANrXwPXk8/YbkxvRpa6Chfl2oCg03/O8m7AF3Sg+Y4MoLij4IdSXp7z41mMzU/T
s4Q/Qjn05hud8mUOth4XjWYHUEw2eErCMdNUaYwCIF4a64/DbWhYuZnTIlT+HRu0
f3H6ZcfYTuVp/5/dJQQHslE7hXBZvnEs8EQqdxqSyxNCOY09LyfRD11BIPIN7m7v
PPNN48yhdcMVt1AN3FMlcwmMbXm2Q6+JXafSgY7Iq2uQ6Qsd7Yv2zIdCaY+m71Y+
IiV/1vkMsxmsU5MHb4r2ZCJ/NTsDzUMwVTcIjlWPHzNpBPj1dxLDllXhy6N9iky0
R/LgToZV+7hHyQElUao/QG4dkvCLyd0s9joCYxF3Ye/xJRJzV2GvPn2oMvg1gECN
3r9pW2oO5QjTy5Pe895XyuHJ7fHm+iAl0AwGxP2+TOTEDib44l1JxqWOuK8kJIAG
BStzTzAwXdeinkZMZtji2CykOHThjDL0JEfsWF782O3AAAe7WWaAR2jmEvd73VZW
7KgBft/1HENMhlTilVubYynMKeNQCCZXhNMr2ZqFvKxQigip4I0xWV5eQWi8Of5R
LwXczGmORuSFeeZqgC68rBWouUf9zYEibgJQmnaOYAA1Le4vCFPkQrfdxR3LGzj/
uutTuoxB+L59YV0nfuDUWA4FLIdkhZYXL5jxbntHOZJEO1IO9DNLRyNNSukjd9vH
8sWMLcvZCE9qSGymy11VfHto/Ec5UgiiNC1R1e9ylzVtObW9kZf+glyKF2b7WxmB
diVZwCZFvjejYI6A81xwtbIvLzsaq13OqtNthtXT3YEwrmyDKeOwwa2C9nJbHON1
eH7jB/ca2+Xxax/KHO00pMKA5f98SaB8m0ka+w3AnU4bGFE0u7VTqliN1+Jfbskx
yFnmaSVXccAY/ErmTADb1QM54tuTAEiZZ4GisGG36Mq1pEePKj8H8/qyjAXmHI1Y
ZraTm8nwhU+LhMgcC2KsZipBDrWZFJ0ivTIH3Y8Alrxf2sUAQq/X0oK+JFnwyqKQ
3dVFmEmDK/pYjZLpPM1Ruojoc6hJ3Rmdp/DZWSzCOiO/4jXgRws4z3p1xYk8rYtA
TTLslv2oyfYNZPAMjeh7b4ymv+iYyS0ZdyFT0YwpPKBSUVtFy5GSwxE7IvuKyA/u
Tbk224YewDgHpwSjv5cjaQkGMTqOqsciBOPX3QCafLKHgldM3QsXzNFpxBDrTs63
aTcfnAyFJfvo/rD3JcCzuxw1+AQogfmLcYKMTdY4jTZ6/sSDwOL+96BQp05bpcRO
7UAiXtG0VPeUVkzEXzBdyNmgZl4iHIy71PhwqOLX8u7yZJedw9vHhG4rrhkOwqXp
MENu/ZHa/Q31vLJZZrmSg6KJ10cwCrzQgjASegjT+kIYcWG+7IqLJSC24DreA7QS
JlrVetPWoW16ani3XgB/VNmTCeCdTMaVAkg2H25IBDYBUeURXaoLG9j1ENtg5Fww
6g5cdxlspO+6R4QkvMeQ3jBHU6th/koit3VDDKS0l60FOrzHojiwZ7W7UPREQnXv
6PT4HmYFO5a6VvYOVrnejGrd6bC79gyztaur2DoM9kcub2IkiuvKNppI/2h+8zRx
2XzaI1Nmawbq5ozHlk9kKK8UkWbbo58jnacVCEpBczFNhD+fPDPD/ZBPGby9dx+p
nXdxS7AaGZC2bpIWE+3YGW+SuQ3whkP6DnZYW8aBuPbjJokCckp3coSdBGHZDY9/
T56aH8lekuVKioZKNUhuSd/mFx2yqsnpEmY7ZbOO1dR0MODzonaVlbslVrE/v73V
Tu0P5d14718hlzeBiaEOxsuO1HFW4D1mb9pSc98lBzpkaXnr/pRghgJCCfk2W6zJ
zRQ6PFwmlGvlzDXXvTt1ejMmlVCMedZFnOPV8Rxd8czoocZab+EDbiDVxSSbUrOU
VYY1bdndKsha6Snn1pW2csIPCvNW0g55NhgkQOHAHDtI83jTHVJjiWPeXh22+iv9
ro/cKAuAfynpGQCesIqXuqlZeiYg85xVinwLsFS1PYZyoR4CUsciBS1BnkLdkbVV
BYYytmoiueA620yuRyzw5uxRzmr78RR8w8r0Zc8ktYBLImvttI5iZdjw5JKjKJGu
Bu0azHTwd00zgs+zYOrHHSNCmpcqx+8C1VidCprRLLq5YnFpiJyD+wIURdFrOygm
Ln2eRmzNKelGWrQlKtudjIkZGC1LehLilzNhxWEWgmMMBAteX/vwC19p6v2tJCcR
828s6J1MtylwDmRcoJRat+16+FtWmpnR0VDs7KklPfHuRoSeRous6FfSVNH/mTNi
14Jy4Xme/TnJXD8MjX19HszXG4pTyWqcaVKz0WVC5h/sbPU5Y4aqIWHBsoTFYADG
PtRPH2MrMWv0xPt8lZmKeEGnVH/lEUOLeDpCaVuxBqrsgmhyHBAP7PkJcBrstm8l
w0eMU4FIzDBBEeX1Gx5+feIWAvCWQuqqMteimRWGx1mfRymSmGLxgRsGMaVsp4QD
Nf/1Asd3m5O0DHKmHCsojbg6UtzIqOrj3bz4bKrjzXZyPMWUIKcISnhMax/tXma0
Uzvx9v79tiLhSxVKzDSOTjzUL0bCSGzkpar1kzppyZ7tbWnPUt9tyWm+BW1eH+/b
XUg7JCJwI+u0q1LJYW4iH3p/UAPuAhDFiiHi7joU9d5tldzLHXQA8t3jtC+nrQEj
LBJlWlcF0jCAQE+pfwoUZMsbqjPgfWvkG0hnW23LP+YAluCdoMTw3NpNkqhbcYju
CmGp+We8TgrZ8v1HON7B6unPJ11yXMdxiqa/3KC+SiOaHlJWEHiMlMoK7bsN+uEv
mTIGwVN0lnZKfGcmXoEnYk0MnSLr/7qCuQ5ftzI96NejDaZQ7v60hjplhs2vK24V
YPMrP6ftZGk/GGI8GfntIwAdnHajh+ffyO2wLONy7PL8PFInQV+/tH7Drerg+Y+2
RVdJP+dr7KE8T3IuL6GC/TnJRdH0yaxZ9C+ll72Tw2PW8nVa20WrOUDxiT+MEQCl
/r0teLoVKpxBDF3f8FrALebwYlWmOz44cQqlxpSDzt6EcYKXat+R9mAU/GMYVggj
KlIZQA0G+prPpaxae147MEmd3wILgZW5M2fs52y2+ZL2ePqwBvRhVxltdj44PAac
DV4B1PWzV6PfxBN6gJ3Qj2kB5n/TI0hrH8fiPzI03gxf2g6B8e8Hi7kRXc5byQXb
H+ylmv1RoGO54J6Q51CjsNz84KeDCLKjkjl8tsvttEm0C3JPQI/pfhk/pjoCATjK
3FVbD0lWSSrFs84xFo4VnGQbfXU0pzVX1yGoPnhREfbPH4hiD/RfDvkNwRUqx+jG
1oZP3sKiAq6daT9RrZcQKWKpKWUhXmzL0inbMNLktXNezbz3ItkNt2Z1NdRc2HjN
f7SsIGv35u4UAhO9b8PRIKEesUU+qv4uzPa5Vt56QXFhjdYddsyoW5zenUW+25Cf
09WPlOFLPxvTfYUVo32oMJD3repzcm68WFVv/mqRCB+a5pkvYdUUg15KH7Rflnny
EQ01hMsGcHAV3K99T7kqOgmZgARaAyLrg9WERFGOMrv8BFmSLxHoMZ5Vc/9KuXK5
Y3eClXf4PcEYkDO45slU704O/4WxFFMECxsk4WcHBjMZMwD8PAsR3PuNPXZ9KFPR
R8tV/GPwYCbsMuUOyab6O6Cb/YAAcB7FFwCt91mYllTLHtXgRLqjt8Vpslj7lZeI
1sEooxDCT0yTUCX9AvSSZHFI4FH+4EmXutpKh9qlvRz6QhaXMfuDEum2T3ob6HhX
ij1kw129fsLzxIyIMcAD2PqHjB4VtpVw7MRqlHYig/pPQRrpOjaAOzQXN2ci3s7y
dhHWRSZMBQDYP3C3lBg9D49ix0Pdgych1x++9ybqb+Bg9M/R5zi22fQRngfBmT27
YzR/aBNnEbXhqnaRuwduvuBbxq+Mg7F7dH6CLsVFzHBT9OZQcRhceXNpPH9pqv2g
iYozpUXJ0ndf9s8UMZif988GyPBAglYxRGjr9YXi3NHp7z0JuJDgkhKfkmhqxklm
RkQ8DHxlVaDmrUke6uZ6b3d23U5MKMH7UEeXvbDTNtQrr9yBoZDUpqVOvUr9ZHsB
cTu9CPzBHf/Hy36tyGOBbbHm1/rgFqYIlDJYSQmPjmT6If0JZiSE9uKRANs2UDHH
hsNRxVqmLXKAYXxaP2a9A5WtCSDHjqqjgIBvC00s12Qtt+AuZGbQjcpldpUnYSvW
IPW3rrjMu9g6EFwNA18Kueg0Siu1to5nSiwnWywSyYG3i1lW/m93WaLF0ZhZaE+z
lz+BVGMdpcmwHq1sbRmStYscMfCGyArpG1AxxSoWJCAD2EhIN63QaSxMfNbFs4r6
YmjclNugKy7decDWvxNfIV34WP7Lowp5LoEMgFVkxol5DbjEh81Uxjcd45IZbmSL
2P3anarGfq5kwcEHhmBYQzf4VNmZJvA/eGs9p6c7Weyso7vyQ9AhC8wIs2Fu9zaa
g2y15RMRDsrk7GaKm7BRb0IW8pOLXPBGhxgphtGPdXZ777A/VEVVW5IXbKr99kua
7WJNa3QV9DYvMQohLd2+InsBWZMXr8LooLMdoIEGi7Er3M3Hxlm+URzgzs1abTL4
SuOmNZWmor5UJi9gwvQMSMvS8pD2hrFYcVNCPbpC0IhA/I9Qv7PdZXFJhH1vlt5O
CzEjWkXbuqYjUDPGWfVO0yknzUv/Kyl5UXTadsjy3C/IAnqPLE1ZxYWklLlTZvNW
1zWUSGLr2uJpqdnHda1ihKasdHRhXzl3KUgI2L1PS6GE2uIVeACekn2IrZN8vOO9
kjBs9UECcDVdenO7P/+Cg1wW6zuYvqnqz1QrDT/qNWt0YKmAzMzGvMULApFq+WXC
53snMRJ5niGk3balS6Oxu8GuKY+OS0m1kSB3yGG8RhnAiZC6F40HVqPszBLt4cUw
Et4vnKYPmrqPC1t0Gw3a0BgODfzVW2R4EahGjwl2ZwfGsk0arRf9YJHM3wNZAToA
8lM73PPhQ+beClZZFrp1L1TnUq58VzRDwCGgbBs6tHWyMYXsDxZJSTyFFZntPGEQ
8VogpCjJNgtGMg3trqvupxmIqsmaBkQJxJUXpvk/8gCJHACbxDnm7IixdT0NPzT/
spHyBKFHPEFKg9ud1ZV9u5Q8xsYjmXgDMu8N560McFBJBVTmx5MKg/EfhU4h61mK
9o/fyilujkoJPQBUoxaPcmU0IPxdLwwk+hnPrzO9GDpVwt6G3hh6/ZgVJZW1Fa38
IEP9lpqasVvf/tk2ptOUJIpW+P0FySlbNH6rd+v4E3s/jz8P5bDxU/Tb58enEMyD
qyqe0IdLfNFBAsw/4Ai6YsDsFwQptcKQuo40Tda8JyEWkgIZXpB0aZxOjxOlDKpC
/wC9SJu6PQxkQFPgKOvbI7hfzVD5KtUWM/FJ+hRbBOSiB7/XQJ23ClG5WtPUnfGs
tgXyZt0Figcd1oUUi19LZrofMiBA3QdWYuRoV6GBHEkKyrPltkKzQ2EMgV+4ytgs
3UhPwo+XJobZ0UlLRF0Xpg8iXgx4zCb4cg7aYuWOmq5r74n5GiAwjRTgCQg5D2ig
vujZ9YuHEt+rHAX5KEZCBJ9T1yi1dsAUhvtWWr2T//6o8nzTF8XuYAleW9dNJQmG
v9qrMIlMR/LBwKbRgwNU7m40X4Gn7A4xTnlydAll9aegR6GKGoYVeoPEVOX5EEfi
qFRVDMT9ep107p+oUyKpaaPhqzY+ofmNRYA7cssV0mHYtqzxsa3YVqi2tNLxAwO2
7dgpnmC/elaCKPxvFzpXf8Y8VHAMegYKM947VJqk1GUHu3IZPhhcoiY/PhTOvt22
VV7lhplm8mvmihecKXo+uBwUJXwdWCOdtNQzoE1/idgzYa+d6HgGmgq9D66uxWln
TdV2YM07zB+hyDNgEM3L16HcoYXgEnGHxWliZJyyebkAXfSDwuTAab2BZf5nNETS
s+fLX218CEBZkaSKyE6rXcVD9MkTH67CrvqdVkF01rWSwrirSvH/jrkcZVIAmUao
pvB9JedslUroUWPQlMQjfYyGvGM2u0M+lYGr2XQXNPdfyse3s76dotC+mMoB8bvJ
R1iptzPd4zhxJpE61UuftjfJT7fiTJvs4LAPTNSaFtd0hLgY6paBjA9hdi4ZaNUa
Kaovk+SpbgunX5nHplBSka+ZlQ2BZkLMI7McIZrYp+IbBuLjNvTHeSZX03L8gfUG
SEfBMaPB4bexrW/Vcazb5T6VltKZV21raeLnFXoyg4gpLacX9uutkFhwf0Ca2YWl
00lOFU8t+DKMVbuLJkpG7Yde3ZmCZ3Q5BtGAEtE3Z0NzsfKMSHZL2aQUy+F/sbuk
QNLIN+xTrq086EdWEWngBMH6GRRKu4O1d5g7Mv9dMYWM9ZuxLJLoezV+tfsfmFVr
tRRUVzq8PM2tyozmF6ssHpxqW5d4Mh09F1Ie5Y35vNKU3qamxzp0DPIKMQU9i41W
rJmtAuU0GSugmTJHLAi5MX4hwvRzgteHX8jzbkD3I9H1tYbnaXhm/3/FMx9tfPQv
ght2IF5W04L1HU/qeZcCjQAHItXp4i0a9IXBlUVlguHZfANZhugtsbv7tv9g7R48
tH8szjtvhUwOc3QpLgG24XBAdw6Q51vfwK1gbdfCeI21dfzDJUCDYlYvM64wMew2
HOPoRwPc9JD59Mbe9sg7cyKEQL/PfNC7zKVuwPSLXzcDDq2klLmRrGrVA3CTXq8k
jYVepf5wSV1gkJUXY01vJ1NZjWxseZvHl8gD8OvN1sl5kKV6tDqSREH9gBX0ZfeV
HAw/6eRBLiauHXavNRFV94gsbgTTBWT42DDa2eLeI00mK0naF4yJ0Nbmgp/Ku7bR
6R4NqTsb1rGQ75J7wCORqzsG/gvD1In4d0iXcedkjIjk19Fyz3mIG6L1eN3Qf1Lp
XFmvURkj4mmm8nacyRhmUGnNShaUos0EPQeJAH8IDCjdza82+Y/XG47gehH1haKP
p7FnKlqq0rbeVZESpac60YP8AEf6E7nSwwUw1opD/jNrP77yeJwlpx8mFdkhcJaY
e0BMIcMdCT3FsuvDDWhITh7WoSWH0aSA+C2a/AqDeiBXfIxYnK0L1fNC2BMGxZgV
eueEWtoOCn8CFL3880uX/DAsRzZVTZXbBA8adExkEKLm6nK+6AWTJZKreeNBEzhL
fwHA4dHoCH4SZCG3wng1kAlFGVQiu26d4Pz79Wt/dTRpDuQXy9keapHHijO+m8TL
2GArHnx9nXXDfYnBbGTcpXl9BS5/kxQadH8ZogxlmEWwBbHJZLrnYZTnJh8Iw3N+
bUy51h3vUhWF5uFw3l6GDCkeIqO5o9D25hSff3eV+t7hLH/s1g+KfJawK3+zydU5
qQ2HzkvE07xoYQmFnXPOtafzDYm6z9YOPxqjtKAkVN2qV/UEIfmXFAFLbBnLFuXz
5eCO/efeYlCK8/Fj8zQ9I12J81/3c2+mRYgOK1Q9CwpsHGKukDtWxMfEmTbaukyf
tUCMJH3aeYwcqXSKi31IT2PshT/8XX4Nd7fmHroaCbuybOLrvkJipNQiS6Lbhgwx
pJETmQFBh6sy0egavDdTlhh9LQWawtwa8e3ZHwwMdjcDrTX2vTsCnkfr796l/eyG
fOEBLcvqhUds/tUDDVFbiBmW5N6uspaBTE0VMkMyo9EwkVqqD9dPpjVP5aeMH2ur
fmw+E2Kq6yZv5dsBnaU+uwlc/7qaGq/jEf9l2WShRJeRi0RByuLAVYercGNtuq1f
tXNmsvdmfgGmo9S8rkn8NQNOhLU1d/8uWQgJL5OK2FUHkoSgKrwT4Rf4Ck/AIJ5+
mU7acWtsHE580ixUFjJKv/O+ZmEBxPOTqy+9YpaQwiQx9Pw6yffN5g6xKXwuTFtQ
dlfac/9fiwRiLNUQ4EveQwK2pgvTNabtjciCWkGoifWRybYq+75BEyfJaMsTKlE5
/fVGTqO4my5Y7LK6aZhx2YwVqPcfn1NehVOA7gU248qsMi85EBicMvOmnNQjLLrz
8zb+mC0UIE+1R68YRgWg/nPi9ThMTxDBHVtoeFeUIyJx4mAZPidAjfDobs8rPJGN
UnZTV0/4hZIMliiED6yozq1tPzGM3laE4605DgKIKvjyZg6Yb6/LrY2caAeB2T9y
5e3nZj2Ek9WCi6SZ0MbHqBm/sAbCYPolPKk3NZpWxscdPKj5IIMgSve9wFkPvmOP
KG3SbMEttIMf4Qx/oRH4CkxgJZQo13s79xrNJBApa6hAEEQrAFjcf4VkVRNNSXaV
A5ZhLA4/jR9gy77AcjuxrWjqBa6NojCyMP6iPrCJ1PJzcbnblBrUSRyKEIpYbSLS
M9+ZLwa9u2t9ns928d4ib7CP4YLL0zqECpdRAiqemCo4r6P3E2XYhnS1u49mkVsR
D0vRPFBMTnxLK2YMFhACIU0hlf2O6bWUx4m0JiKwwGrQPP1PakHRcO7aTx7a0nHh
2sxOw31feGEfYzwXpgnMzStJaBRSgi14L20ayjEhvy22XsIq3rMzQLFU9bU7KjUT
ZJsN3eVuS59vZMZhsyEAfWYbXbO6T32zPlwUbzUx/yQ11sw33dCYnnRaP1JEHQwt
LQ+Z2x6lK2ReDeu8CHkKUTeRKCRerTPVl87q34MBES41qK+aG38mHMtvBLgzJqut
sFgZVAu1pG1IS9bfVA6C3uAW7F51fSkqYszvPmwhY+e1/963HUL86uzNpstbEgaO
mBEJgNAWf9KKsf3VZmCFyrqoIC3+jHXI8B2ZEisWZg/RsMpVjDnApLkC870HsAWC
oltiegsCGK7UCG3WZH6KN0HIGXtyTCn0hyaG2sDvOU7yIFQoGWQvRJJJxduSEY1n
zfY4sPOBa7ZfoA0kLKqAUtT/lYYSnKLuf/lInWTCgka+1KrkbX0zCVPjfngS0u5w
LfDYSFmiVlwMZNdQpmchBe1mbsGW64izxQzZ4ARnOvlnojRBBD1TTcr6MyA47k47
x06A2eNq0mafsMol7yhH4sw/ltx0kQiPDdQlyVSH+Nw14s/unUbvDTXyp2Q8iwF5
sZOjUWK7prd2VGEpIbg8PflB54t1XNuhUcw9/Jr+BCfhgmA0PJSgTIOD3vwg4y+N
dNq/fFycviwVJyoERhqWmOVdM4c17mUbN6JbqnNNHvOfAXZCB1TGul76oCsfjD1C
5rvcBvrJ9GlKRlD031jxjln5OK19vQB85rKF259kkr8GBe2CBuDsqLWNNcGMhXnR
YBg5rXFVvnhvU53mQ8nao8Q2RZsAbuKEPjawpXrW80+aGNoJG8/leXR9e8FJo52z
f6R3XccCuzaUWZiNM9Ni/3txLyHe0x7QeOOd0A57fDRvnc7RV8QAh9wmEpIutHoY
spIqAkNILyitPehwGFGaeE7PcZj3CV1MuOy1bJ5A8hUujnOw4+uPzIeeOEiwtDr0
OkIz/JxJZmCiHjzbjGLDx4SU1ZDjambfgObEMKNznhGyBPLCJkZSPBZ+JHvCLVlI
b4JkS/SrO+i6smmKm3/VTk+RTdXqf6xITi8k3tkGkWAA31uE5Q05i/p2oyHZ7lok
j6+qGmU/FnmbQfr12mgzL+jaoHyY+Igyjn4R+krxNS4Hd6I4nxiu9RBrGJGeVEnI
bqqpEnJj+kfsKUUNrotxSIA8dBKyjDm2G0KbWPvGZm09J5UCUed2RejTQ59tUWZZ
dZjsekvp0tV8x8JKR3Ita/z1FzbWruqgm1iFBr3mJDQZR+zhuT41cvrp+6Rws9NG
ZtWIfqxgo9Cl863QVsn8nZ2et44JzOCErLAMUOTvEWiReMnILR/s3Ks2Aru795j6
faU+715IPc4E0jVQ7PLv2fz/88RoNUFRPhaWnGQIV+e3YzO+c30+/fxaMdSyxHp/
6aVj5K8/Z3pYt5FTTnwP7+PaR7DnLwGztqvju/peqsmNWjCPJOjeFDc9Ij0YMR4p
mES0z2UiVoO6UBhkZOtJEisNbM9k5R5hm490NaJKeZgizOi0ExDpnVUVCP98Hfd4
jFbXgyy7OWLYB3dTeTpRx3WbBlr0JHsVYygEaL1wQ2gvdzNXnHjSy3YG/RhM5mDi
39DbYvwEteyzjAu1iEwltLVJFpgRDKG6mfWYpHlBctbV0aesb4fCLN62VSez0xxb
wUxWSvn4heMuyfZllyXLLmm8zCGvihQZNtO71mXMSSTd37U5Euhwrr6kGI1/u1CQ
gdM3uwTW1KfB3VHdKSA/ZsyJk1IGBxWqhzYJ5o666VX4aS2E/j9RV4B8IM8rSv25
LV6Sw24xraCdTMXBaF/qyeQZI0MnkzuNNhdqMOShwsXxZoXmZfvEz8P0LU+C+5JY
8TFiNk0URZ0icgj3plPjGjHAZClpRD43sg6fTkUaqkc6r9lyAt6pDFm7Xd77R0kB
EdYexhuKzlYpmuOPmUFI+Y8qgBClG373HFWqQQ3cuGfBfF4+2pISTIo3RHmgVfr0
gjJT7SbMfOjn/6aGGOVVsvuleOTQFvYFBeTGeb1WagmnUQ1ZZkcW0PT12GL4vP86
bb5J3ucIg+53SFPtDqHBqv7lnn/Yq3+R7JLSr+FrZ2TEZAwcsOtPoomuLH3tkNnx
DA2Hgg25MmPOklG9s2vD7q3rDF9pL7wRlT+2lkHB5xtgMEocMJQITFENfNckOr2D
sIg0OwAh4LQpphz4ozfqVC61ByhnUVYMqHBnSMkK55qU/D7JsiOLdTXxqVbWv80Y
9+sF25bQeC2AtTG3HMy+0+AuvUTqMYrQjyjZvSwmvzOxXbdev+OOWpuz4+6NQuO6
y7d6MfZLtBHXTkxMA+bSwo5jCoZmmzF3MwtgBGEQJvlfrDgQPIEfH9/jmVXRncat
hnhRDIxSvMscDbHld5597wk4OxnPhusKK9W3+0ek0X0td0cxmGRJP3l/TwivqO/R
/I6mFVcp2A4Zjeye+gQgv2UpkoFheQVD7Hto5nV4aSX5OFV5fGiwgxOTN01eAOju
Eosrd2Zq3hz6GbPnANP9etMZ3yKX3xAC8J75HqisVv2A03n63k0rfs8HixYVHA1Q
zfb6AHWA9/TDpHV/watkvz8v2XJ2o0W+NLzXna7x6yOSsem+n1eFomCYbr4rnPME
dglu57+sbXPw6pyQiNPxXqD7MBgUviCUukC1U3oXBEvPi3RrVn5CHviFE5qeD/rX
c0bbosT3Z6NGw/ZcT8GZOFkx9d9xJs/HOZ1PIXYDjpbuAJhyJCGrFK5nC8yy8fTB
eT78X7BjlEZf0gPTjolu7fEoSR/jZaUckkTbzfHI7MBZo5RfZHoZUx1VFH9aK4ak
ipxPAB+cLQZCKmeu5/7+2RPUYVnSF1x6Wt6hZ3DKmL/vR0+ks+lKKyVx2pdr7+P4
xF26M0NDW8PJpzr1sKkOwYnnM10S6c9z/qCatRlkBofP4aGEvPyv1Nl+epHz4nJF
bPzYgg8/0PetvT6KpaVv3qYFfUB762YzX0dkDU8zKqHQ6KN4CUPmGBVVCQ4l3gVv
owO+MaEAdWTN5tMPLAgGrkQ2vnKlmDEzN/vWvqcfdSjAZ9rZhWMXYs3s/hJTo4gt
vqtt0BypD3tsjBFhJGfNfnn9ZKctUn57P76U5a4xlzbkiPsdqlUt4XBwks4XNip5
Z6rEV7ouOlgTRMuCIyVEweImqwra4vpiZnOoD45kXheEiD9VZKWEI6DW7gwiAOP9
KCaq+DoJwBK99iW/hUhKBJ5aPzs1pPARx7dbyWXaneJ4nkVZLeCtPMOGOP0wedyl
HtaqYTU01sJjKfwLmg1gyjsKMIoNIihTeW7hyltJNZse2KnxzwR6Jb6PBAiledXz
M1mZYEbL1psqHxmjF3VDNjD9UPEZYlT0x/JcJ68IcIvHmc7XXH8nIOuWyCEQZHbR
Su98bKxS+SIN4kPRIsPoIUah6EHD3Ku2dTmUCZcY1sRmEQye01nQLZ3BtKnV++9K
lIqSFuTlEiCJHS6LGQCfes00SSnZiooaonPTl27NGZu6C0/Jkn8z4Tkr5ynI06kJ
Zr6v6eszofXiLP1elrLbgQz36ggss1IlBGr0/0rxWXZJdLR7R0WNRn7htNj4vZgR
IEX3u3TsHbj3XCl+iA+N5eu2IlBWeFdlxz8avdsPU7Zi0dcmZx/x3cgLy9N+UvIc
QiDvv1YgXHMutX1j+RvyL5cMArGfX0CzxFuYrhzuZ9+4/lmtObm6+62JaEjz4W8a
KZX5xMaqLCNAHxVhvqbTmuFhyGLDdTuoMqUIwug7fXfwZTgPqv51a9GgjaBBOyT9
/6a8Gj3bcYmClFGO2Q8VGgTJkDdbRoTEfHPYMv8RFkTlfCKvwGHNEawvuMLnPEBp
FF+9sIngz7hD9sloxh6bz0qXbGeakzF/M6vPwwjsquI7a80H/jwTajTzCoWzrv7L
a8khoJ61v3l1BkQQKCRNfVdjPv2BqUhKwVkvxq8VhbwFi4BrPa6U8NRa+zeG8SSI
4Flu9Z6yVhqUbqsyjx1gl3MlCPt+crpQbkpp+4D0kSNhke3ELUNwzNyXo8mDUD30
uLOZm4LszrmP7n1/NyJRarJnyV+y8TRCF6Xn5rXop1o8Y4PSVOUYjVoyNzvZ6Y6V
3VCVEG5fRArrjQdI5haiYedjRltj0gleh3Zoq236MXdVpbypdtYZpB5fc4QHsX7C
FkKj494asxSsWvalgAxeivbX2a1fvRCjE2dJpfpEUCjxEEnXUyZ6/pvBDYpQygrh
bdyJRuKalHN4MqkILil1YHZlwe51fuMWSdpOaVj4rqudzf/GOPw9VDoXYzyDdzSb
2rbDsIy7FFRP4oBH+6DzHozR/pys63gCOay8J+84xKV3DKgkpq1gYW5/Gg01q0/v
wck7NI5ollBZOtNAVSKeJIC1/lISfn+sXMsZnwOsYbhVh0cl0ju2fsjnV3G0XhHt
ewB6UA1HIs3igKugjHMkb7KX9tYNoZ1NGS8FyuQqRVbYDDLuyg9S54S041TklAgK
MqPr0QYhR5EYBYYqq2cQQqKieZe/4wYQ/JtPCIn7vp3L0cBIY1NPr8W7URpFq+KL
CUjwFQzGzFvKhcNEG9y6btnduwtu1exdlChXNk9CxEsReveQosGMe0jumItU7p80
heS0xn02Rv/UoANmzIE/VUzYNWuaEhufCIxl6jI0gVC0X5KL1DaEp7zRSVBYRxsc
szfw26KXYswniMUGTYdmKyh9J9GukcdLAbUlXIHsriWcm++8kPW/4T46OS/0WyGp
b8PwNtW55YIRKVSmjMuIgX6hVSBHlkSMFoWXedRpKRJWC08RutdqfGCQNkRS3IO+
I2mh8yQMIhh0RumxCvnFzMUKfC6A1KBNvwfSZHmx6Ex+YIJebhkWznCroHE6SzVF
QoL6y+I4MApoWhGWvRQkA2y2Y54FVIwbJlf+LdC9jWL0xLoRhE9MIK1YMPLvjDGz
agN1hBTDMdbs86k5a2xVh5HLen5U9hUWYwsEdcm5d7zSkpulguIXSEFZTlXqfVCJ
v5e5gxlPsQzGXl/H3BQL8wAeasNTwUuspjt9zA8w49EbWKZWpeoVTAw4fJnGLCN8
prQPeBPdWFsTcUikTavCkJQui61IMOborh44AZNHzPUsRATCshh/ULdmoSX23Wcf
7xDYcQyZ6L8qND/oFENcjNDTJ8n9yzTOymLh/aspIlFndEs5moEz5STUFmvDAMVM
bFv2F0A76C+1IUp78A+GPYyCYBd1dWGk7PSgCkgpYezHx9CNgWSwtqs8wBSh0frJ
5JgM6eYaWfRot2DFnJPc8uJIVeNe7fpLKq4CeUWF/sohVeDV+Oh4i+3ADNRYBu+9
nS1l3neO4QzvKDQPKrioVKGBRZQvrzZgWXDXiJ0bJIQpvtAJdrqOOvqFenmQF4ws
a+M1UoV76jwilrDrDMZXGUlc5aAY4dUJqc/66kxNe9MFO4fI0tr3efUO4N7H7bQa
DaxR7LbxSV9ogtv82lFAekGP/0F3FIreOwsdSVYrQ0RqKZfjxExmUWjWbEMnwcJp
SUeSFzKoI3L9wa4Kp+pvBE1b6zkITsKB+yQDZUWaz30UANSHgPTl0BAe2n0E8aQn
u0pxT4LX3/lN1Ovgn7c1c5H/NVbBaygDqOfUlDkbAqVP7E/Hvie7J9hIpjBUVZs/
NrZrIl76Rgvb7MjRS+t6AJkmza0YK5c6wZR3ApFD6E8dh6aWjPSzsyviGlA/cvSO
hPR1M61Tc8ChvIeDIvoo733sDVd83Wr60fjWDHKPkyyx5xnOUqjFmBxaaWhNS0Vy
sXpJ9C24TdsjAhxugdDfgb36eG/gH4TmSsCIGb8X3AvcAJzstsT3rn38gxW2FojY
JIHpa1Phf6rxDhOt6JpRobe5SOa9PBgkdydNJ5upjL+AeCv0YJOMkbib2EBTz4xu
W1NGgh4kXfJh0c/YLb61IFkTQ2tKDn5oICAp8ULhF8QeJZd3xr+1tx+ZVH9WmvIy
TRCP8jMAJ/MNvf24IIv+Sgf9wV/UHg3fcsF/ko4c/jxccv8lOOB9i18se8H0BvEC
q+IvGXulLC4zCMmz7v5ul0RPUSug42g9oRr/MOGKd1mms5maGbYwwlGN1gN4uHzB
LDdcaBkRymvRJcZlz8nvqpHHQ/O00Vjay7tuDRqG8yns1r17FDi/3QGWgxkFoWFs
1ZOEIz36HjqefG4UOTdPCpFWqY/pzgNckQz63R2gTZFIpJBursViKSWIU6M23u0W
a/vb8VxfWXZsiedFkaeiMTUW475ZneururZp+uHD6rx3uifKCvWc7qH98ultJBCQ
8SaqoIF1+y5pnmXoN5CcTViKCOADWRl7Ej3HIBunM4BuXZhNP/hdHKKJq1ssR7Jo
uBCVIOsR2WTeovXKqH9g66tcskYpoS0zTdhjha0e8Gl+PhZm4o3YpsZQPtTtthqG
uELt0R6CR9QGRGPJ4JGg38rleLKcFpXiynlSZLWKIPvYq10gyk+YBSax1jSqRCHn
/RE34xR7Byr+aThsWJFn1sNIgrsqM4pPXnrN4JHd/Ebsl9N7CA6jjRKLB0/hHCJS
AoaOyt/sDU1QugKcMfAAV0E4lYBySvlLHGZPIhy8Hn5g/HqIvP9dSqx7w61jQcGp
Za2enhr5L2NBBpThHKl4YDTpXuBTRLBvqdyC74I3sTfsqKrM7k8qCrp+3Lub7qeW
St8l2R6t2lmEG1avbxUuovbNur8neRpOJIO8aLUxvArEmKC5OFPejmvwsmvRfJCH
1htI0I5FA+W+tnCklxUOCSx82Fja9SwZp6SgIX7gZYbOqCrA/H3pIKgJaATr+Haj
MimPLNtkxrZ/6G3CnYyiGxX5ND6SksqrQXUNTaweIlBRnoIber1T/jEGeH3j4hdy
Uk7rsAl/IDykVBv6v7wH/jxs7Bva5xKAvlmr+GcaI9NPQWobnoY4svblT7hyxvbx
ahttYgvW1h8J9TBU1/Yi33GlD052dMrl4aOALtLmRZv459TcujTuH4xXo13Y198H
2e2J/mFoAk6KK6Zg2of+N1K2uTbQz887ZzNCkX62aeiYkxLu0Qvw5Wq0komI4L9z
8rCTDmElVggI7JkRXMpJKiLAYsaMITO/nWVBYNpejHg/N5BS3FKNYnG08nRoR2g3
7IRJYfDcMEfzR5kOG3abAZRXI3U7WqDRKV21GT2Yt8gBeGMIviTPjSoBDLlshaFO
GXjfEtqRKic/YUVYosu6oJd8O8SF9MYptr7yZaY91k9Nnul7PRSqLq018VOlqwz5
X0GDrWIi9nCVN09HyK/ZmE8KQ2SiuQR49NZyZS/ijzGM3gDjeVJ0a+OQejuUNfH0
radTbPlCAUIhvWtal6oKN4m/0L3/UFtFdcAj4Uznt1+4cTJOdlxUNQH1c2e++8Z9
eSD/Fx+ZqE3t2uLwWskGBuHdc6oObZI+y8wvH1729n0p+JlRQPGt6iaNLOYyIAuy
zcR7m6ogopF/vKTY91tq0G99/YZU3JUzB9iIS7yB4MOB44iLi1L4nXg0Z15JYmK+
JfoOvPjmUHxblyzwr8GcUfYwi1SRxQTmLCcVqhgZiCR5ZjQPa13FAkQii3r5sAvs
j/S77vATDAocL58PSzSxUVhttc4wXBHCZZnf0qW4iF47TEjhKFdqgBQht+YaamJi
Rbhi1MAjtw9XT5h5B5+KlKoCkAQtT0wKvE8UozU2emGwNnI/E6FewCPkZKPXL4AB
cNzSIAMtDPv8ML3StWooixyRThf+ssqhpxunsX3dC5z16iocSd6Cq/U3HYItFhD8
nyuvPE/Uivv8pi1jn26SlaTIYWKQ69QddaSk9lqIY6I8yZypZ2L3l+2hlNYJAXa0
Vc3GTcNc8vp5Bz7BvLMfDi+Eft1Ljmimjwh8K1BCmLebhu2wBSnShLz4Q+51OFd8
Fym5bjp1Ewp76JMG3PBAmKaWRmSTePtVusSlCO8GuGTFJCM9e+7eyK9sFspXcAgU
4mC8iceVCNeXcCAVwa4Gu+oMoeZeIAbDeM67qTKZna59MC7Jfo/+DX8LlZQVI99z
676b0dnXQSTUhJMHhJTVjrIP0CEnLN+yABHcdD2YVzsG5+Xf5QHf6sXtP1TqR/Ig
I4QNd8gppKSLYcukbptq0NVf1I0PqdLBjNKAbWqSqkdB23v6+ynvCgIqcygX8FJa
eu+7nTmwcgxLgZV6lKjvWiAReALTu4+4S2sKdndfc8vftdYs5ry/3FBnpXV5y7u3
Fs4plSqQAueARPLzhTJeqaN3wLIlxnlxWnJeDZBma1ekT8wg5jBgid8FrMn3ZfdG
oJpqRkeLw2agNSWjlBQ9tgdB4sTNUMaNJ+mri0oCXjscqKdg0biVUcdG+gKeU1Fz
xkpnKGP/n/RCX1IeObz2QYgx/vLQND3EMX0vsh55I2dWle2gJAzzDY+Gku51vnXY
TPtTLOze3hDHCT1tD22F2YSuJ3naDzOihI7hnZGgRPyQCcQQ7Q4Yr+reswEV/7yG
zldsF9uerwgZsaSw/7sbskkfBkKatvQho5xa0FaqZePvaSWBC9N/YJWBe8Ak5YGe
UOTVSDPs1vaHCBmDKO9o4kMiOlDTVlh0B3Slqt4pgiUYRSsqT8bIVIdDcjwic21x
WBA0GrMNNkyvYSlVf++fLOVp3fH9cn7WJS/bD4DmopyXIQ9ytRBYlKauEVudh0o+
FQfXx1mwYgQRaAkGxv8eQVJx5cYS7+DXlVe7D6dp/PqO9Z6we8jOdq2ntWg1UP1r
+qJqgIQM9D5dvDvzL0NS29/tAranc6UXWzLyQYFjHQc4t6jsnTdg3Y11DNIrwHb3
5DmjcQJLci5fc7MoRRiiVkDQmYl0AsjYHVipGzZR+z1gRrlo5Z0OPqc5WoK8Cxt4
SP5yjszOrVVvzrDUsronTcVOsdn6f+GoKF5+wDbdZy5oTAqrOePpItYZMHtpZmQI
S1YQC51/6MvOL7A0rR09f8hZf6DmAP1iPEw671QeOeNyIuVYlVLuMBbVoVjPQG0/
hpGl+KU2kiqq5ZV6eLckoEb7DO0xcn6qgNZxIKokLfHmqpRIoWTxuxGckS/Ky0Xf
1otCLEuTwnT5UW01lr9pMZz2b+q0M7xG/cx1RJjIqGGvJQo1TEt9uWwCzeOpmXr8
oMc56/8J8rgi2hyP9yPqOUUawpQma3o8tL4xSObVfEi+hEeoFwGvTH34Zwc8pkD4
bvdTQ/qaXA4gSkPx1hgssqGXVPDjgyYi612kNzupglmhMQYGBfD2C4iQkGAEedkl
wANEsVM8oawMLXBWaBEOnxeqdYcV3VtClr9/zsA9+stoLpXTGShPXfh31do2ADSg
mjYmaq/z4M3CJKqmmUJmCzELuZ7sHwPpnTILRrd6esiP5MGrlgnn75Zo9SbCcuk2
lvovHVFKt9SeYEBHil7BGfakPw+EEvfRDt/a7N69e6z4BSx2gjG4ZSJxe04tfO6h
tc8cSno5q1Q7YHKSO2tX5vaZ9tmAjFmSSKMNWdHL/HuzAvztLneIy/I0zO2Ozs+f
BEdvI/XRBbvfcU4B0MAqOg/RXkbitu7peoLdOaDICCgypZO9q86Ebug7qeDPJcrQ
p4rgthpESyqbE2x0TR2m4UxdsTXV6R0EcrHbH61bb32E9xHm3Uac6UEIyLCqm30n
EnpcuZEQWw0U/Q8P50NQSpHrC3FrqxTDrs30BD4KJuac8vskfhRA/rr+dF3D9SZr
HfZz+2MgZA2j/VCk67I5PyLeFUf0KWC6HBztF1RteeMU8PtPqNICMSHByGUWampI
TZ+ZjY0GiClA9rhtJ++M/rmKX/fYFjH9LRzLE8g/PXc/YlhmiGBIVfu6Sq7ihl37
FnpJHPsFdcAVWKmR3aigpOs4yyDHOIDEWq9m/VLH0jjNwjALuByTc/dwvxK0w66j
u5EOjxmjEpNvvwem0NtGTN3Jn0k06ZABIPO+Mi6Xwn24fz1xwPoNbdrsx3GJMRxU
T/dXyiZQIidWd1L1gMQgaLrOZBk2ExLaFD11fOWCBa7H5YKd4CIvvyUl3vwozCaS
K0M87MOxhya6+4aZlgo9dvusElzctsH9WEkWWymfQnxKR9DrqbYjDiL3MhW1XLdZ
y99XL5aMlySkU3sWsq5MoZrH3q8Llh+zUm0guKv/SG6cKkQbcpSrVUO2zfzotUVc
q1XrA7Q1msmAi1vo3GY9gbduKGRatGDQBLbmNh+mM7n7CGquUMMf7bdEzFnnUctq
PAqU92S7lvf5kLEmzg55nZaFS4Zhw7pyA6imiakf+Wgpd1W60Yn3jFW5RaMsgC6d
WeUC6JlZ+hKapKXjmsxb+Me+ku9UTH8DRx13XzqZGDvfNg9tqyldSBeL1tnEAQYm
uxxtpidXyr8xF/emjpZQrWKP1itcqOfalPZyEBNiJfcsWLCnDGZn/Deeg4pr6zel
h2wz923H/EBqLLQzX5ierbw2n/hYVMaCKsAR//7xlGmpqsUOUdEZm1UbpuuVzjWF
B2ItO/72b8nie6btTwlOKkeRDw970fjoS116zofqdsy+EAqaPsHjPJ+DHolrURAC
7gol43KjEWYUe5Rg9bltKEwAvdeTxEfpbvENKa+v6YPQP8qRsV2aIUbEFR/LBXiM
/WKYIGu9OJU6Hl+pBJQMu2SQL118+0oxn5S6qwKH7kTDrYYa+YdGYv15ufZ4EF4R
ZcRxjB9OecEY4DTLQYyuSy7S9myOIeqQ7R1y4mYwH09ydav2NDJqcMrzsGZp9k5o
dSrXqNgndwBGUw0x7ek6J6g+9fAe2Tc4ZphfzhkfMACVMYkUogEWLgbm+54vUWFk
2jWoDkjx23+EhnJ4aAoG4Ga2bFKVFMOPbGTUSYNrrBl6PgRbablgLzbNYImCwcJx
lP05BuG76ApzCJBS4yzQBdlaTsCXA9mhEoJWtfUQ6N3z4V5luIb9uzRwWDV3OzzP
JbgRh7rwZbld8ts8wC4EDwdjZ/mYlu6O9sxcPJL9qpGmM4rmBz1dMt8uV6XFAlTs
9kms3Lg5L7BmgmiC017Mm9Es6/rQ3Y3iRozockUe1sO7pFaejmUcWygwC9sUskox
NI991BnJfa6DzLt4wn5ITHQ4oDKFCeg0XWOk2cgntlkCvGFWMvP2ovp6JZpHk+Mw
Jqdq7KHY47VTj1Rv9GOuGLdjhAOD0nTjfi4hTuqRsu8yleqijBv6EDWNvFwcyoeT
ChuSxRfCESzA/9hpkYmJ/O6pwDGjrVGPs4UfZAl+ZGw9QbGkgYizsQ/BuCiqwVpj
Q/wVUoL5PfcBKG1wEvK3opZN0il4IYSaCX6ZDWWE/WILCvhN1mPW/otDx/f6d/GI
fGVVSqD83BLJtvoeAOWat/q0f9Yjq6lG/4zhZ8JScGK8mCN9rXiyBcwvJEZS+A3L
f01iktrVUQycqKg2wXBiYMBRvInliPtdgtf7tJ/OssmqYY8/NFPLUtNECBenrO/n
Yei61FRu8pVCBsjZm0r9XqT7uUz/saiDxfwnJ3zrPygUh1acXVKHBh6HaxXZd9eP
t/rIuF4/hH+TwJw0+0cM8/AdlQfT+Oqn0WX4WV+F1Cvhg7MFgO7XIdyji+pE1PsX
JBuPIfSUBdM/+ESi3LxIKZ7gzMoRnuLo9mewGSbGIS/9Lze3iOgdB1MnTRCK4MwR
7r3qixt3UyWrlpmDtdnXHQQRlLGJvTTa1aSUBaLAO/GySv7km8ig99aJw9IFvGT0
0oGLfExKPHDV4N8ZzFXHcF+Ohmf9nuDmzTq5g9U+4wBSVXt4FT6A6YwTdkWVNx7Z
53KAHmozfNhm2rsgOjyC4LNQpvr7g9rDJdzRB8vqmsERY5SWSsoFg3P7dRS6a9Lg
QgmF/kdJmOenDa8/ar0CItqD9jumvjYgGzYDVvfonDss2iu/nM1jI1ykKnCxL6qF
pIbWPoKT33kKNK1k0SQnjuYnzaCVGMJXpBYmQrYllU6CI9r13PFpJptMWDAYk0g3
0f4fO6B5TnkGZyb8NPFqM2+UZam4ZH6RzSnb/s3CtVQd7oAIl2dnKkQIsYHnSMjg
NtkYTpprXqz81P6fWEQi5oZ1Q9/xh7gkoGslMF561i7cdQ4rvxT/bzM5h87WGxSe
y4ENtRikFbjGF43Ha71wqKBiNZcZZozBYBBGkI53xrVFprfxcnk1UZYHD/d3gFp2
yA6Qby4Ok2TzC73vB3VfepvWuxgVoKZT12cug+JFU1bcQJGDfi9fV9DJEZJCBOuf
D1irgB6esx0aq4Pj2a3mLeHkiEsY7nocS2U+MCK1AeSisxxXDYDEbacyMRiSpx4q
ZCBT9NbEoLsCLeTGewOFRrg9x/OFcRpmMul4NcyKoJ1t6ga6FguWnS2mmljvluZK
+z7oB5kmZPDxpUEN4I3zlbCdZ0oUhK8FJtoRNmJiYNDA91rOBxorvUbXEXRZZrNK
YQa2c6QBV4MzXkMTEg6/sNLiouY7I5491mXWTmSKHLxGMy/XM1ctL3sJuqnOaAYU
Z5YdX4VqH0DpHrp8fzlfgZk1eg+3KC2QxhyNuss27+6mJO7vNcAmvcY/wgNUY4SH
8SzQzcevmcDei+00V/eSpQNS054cSt9oh+ds57ECSh7IwNlYQlXN3OnglhgD2jTN
vE9WnCsRxKZ4Em4DRdjCPUcbEibZVAgCzpuWQrvC2zddZm2tjLq8lK+snTQipJuN
uJYuEH6/mb4EPnGCBkfQLs/mD25Vow5ypBYrTdkuYUryLmrXjXt48/Q27BCsAVE4
E01JOtpoIfMRNVF5jAqgB1VCANvtwjiCQeMh6qJRg/JFKHcDFqagbbcVAB8ouEt9
KRT0psb4jPEYP4+fIyec9Ywt3MwTlVedmuxvQt/ioOPRlgEu2jE/p9x4WBXzayja
hUA2oYf9SE9t95WJtstaG9v6rvRQUNjTYRwwZc/1Mi05hVG+ctKVHjkpQkD6w2bb
N/1mvsro3belFAbJtoK14Lh2UlSrkbu9XxKGxrOaSRuemUxa/jzdQVOCH0bfRZ02
F73c0eJluf2kbLpKsd/YoHdWXpBT5PvhvlvIB3MsEJOpeJ0iRvXjyF3zDNkZTlAV
/E+ixL+fl+1smZACYWvbb+XSKOcuRNQnLClqYNzDH5irYKzmzsWPYqP3UkOZlryO
hnMIOxXymS6eb7LwYvxW3Me2BieWaqE8sD2BKJOwuWfbGmTky1hJ2EhD+B3GXg55
m34JA/9gDzFZxDAec7yRxrX0cPVJAxVhWZivQAoaIA2rL2KO1H7WbNbPFdeSN5T0
P6Teqz9lyOxHJqjCXbGuaYxekkw1uHD8HnlBQPmzXkSGGCwvV6REMQzzMT8otEpn
APdcjQedGjCtRQmh3TSNcl6an8M5IGPeZYLNtaeb1lFOsp1urYmOn5CQxOM4MaTQ
KR47WSGp90YhFeo7OX7JNdtPmxxl0/+fltXxkCYakbVSP4Mhq04e+E7pTGGn8GFg
vThtWPJ9LeOoZj5CVSMz3Uo5REYzRfQPvvi9BRFbiyhGMWHIjP+dFJwSZCOIOe0n
zeYMOmlQ3pWeE5UW10yUYec9MYGSChbei8GZPYEeuTQfY25z0bLRnnP7cFf5eqmL
mVCUfvwQ2oZLaDxLYvzekMwUSrDN0n5A6fKYD999iN+5r+azxY4TDTE3IZyCYI6b
B5SPS1HLB2wEOr3YGPGgXL0LuqbU7FIn7y3jXfXzVyPt2/gHJ7Ax14qke6Qc9MLW
sdMzOh+iJqvCxCghZQhtSDWCUg8VBkd56DoKI1g3OTmk7aZP/dP7bF7BZI5hVT0i
6EBEmpt03VsmyCRE+g1Nd+30wkUi3+/vOMo2oYNIEVEim4L5o+ebythNoUsPZgNX
c37iNrSHwaIA70q5CmtCdxV37uJ44RwQS/CP0FzNjui0iA18pNFAMOmvVmC3/pHj
z2U6Zwm6OZ7rQqU4MMcNYOLyo7UzLRCrGtec55LFWJcr5DNJ6IlZ0meWoJffc7c5
JJJKDBoMAQs97vEUUM7S5i/AkHSgSfFp+WzFlq6PFLobQmk8qtIOPyZpkFkiLFEb
bJVoWBCPlF4dktZvHfaFx/2pPjgc+l2GSDXmh9aYkbZxXxQ7YL1UfEPiGdII0U2j
F7Gai78y9JrzYn7VN4pnHRLhhMSQxIegcNQwLaXuaJ7vZ9F7goFQ0uMYmDX1TQVr
X9li3ojF0NgfwJmd8BhWHD5ALuuSWi72bW0XER2rxMPGzgGNJ/UF1Z6oahNetG5j
ie2Hj4iuMD+hRfjGtCKrP9s65eXZ75Iz4AxGp0lQ0P7dwi2k2x+Aj2art67cjnKp
tojIql/chDfhhVSERBQi4o5Y/VrIlC0cZ9Kkq08vztHOZwVgQAic6v+ToGzfGd79
zGj71vnM2vXoftS0ZyqhTlilbsnxxVlm8pAfOLTU5IGNRA8urpiCxlKvWMH1HYRd
mQYztj7yTxr6AA6+5TwpgftGAfYk3Z2SFCOH6NLEeLTj6jtM4mrfq3KDUXX0z8x8
+ffSyB3VSlOS5OVxcwteEwpxf4dxnTUQoaneYCfuN9iKIzgx4C30dmix92tBrFWB
utXZ3T+NqIJyMV/I9a7BwbRAXByhmplPNpMPP1AsBKvJWKzdc01HQ0N8qfgRSbUw
QWqbZLRZgbhLNU4Ip+Gh92mfBoc50MBdfDy8Xj3cuMAPapgRHkeiztR9SRjbkOSd
4oZ8vYhXTlgk1w/7jfDvRb0CfAiFq1GYjYLZWaSnnTdfRe/bsLXzVKjMZSBAf/07
9+/G5TsefUMslf7OzNuz8yL4FjURUq2monFWZAmlFd5P5UHgKB8Dvr9E0+WZ1oFK
i/exoMOVAaalrTFBcUy2N7Uwr7WK96yMa39+ycSbhUNr13zD8/gGSYJm0GswfH70
0qqrS62UPEK+xdDQTdNzFm6lvvu0s1ujshIL0CK2u2oF3ezRWr0ZBIu3VBFY3CVV
HZkApw+OrffaTZTB8vtJMza8jBnw4b4kUTMxier11E34oWGAL980Ub+aoWPMrYhw
XYesIx+6tNgle6Li2lCbRRSLS0tXx/8UBuoeGSNT9RXDUaWHeEZEghZ9cEoO7Jeu
xIQrWnB90mlo4Ne1blOs9CAGzopminVhPzTKQdsxvk0deusgSDjwXsNBWuqkIK6M
QbJsAZ5C+2PAZjNk2XjH1rWwVV4is9KkO/q1l3D+PagxdezSoKesOEKomXItYz4b
b9LrJUwdGhqVHiJtubiZxe1seQKxuMO3c+Kx28DTu505Jyb+KMm0Ya+DGRrtriZE
gzdgMKbBBwuJ++Q67SeGw/Gz/THgkko9/xTzxbIyTPe29zSNcdLxHSBvtE+DC35Z
D8d1BejFg31+R0E1VsDIJtjxWy0RsUP4YPjA/hcXhK9J+STx+c8T0KRy/IVO751I
QUFnRIBwQZNSUaHS0va7KQ749ddxv9aq+AqxFW+Recssgb+X0u658j/3qA9mt7Hf
kzbRnjwCEyRZPOluo4Jb/PQTtJ2/QnVS/0VTueAFmF3HoHG4oMlIvlh9ZHCih2ht
HMjgYma8tkDRz3S2dNyU8zoIrp2j0UKm0x8gHxQYdBGjfyW9XBtcELXToC2RQJ9L
Kt3z16eEOoaRhfCkjH2mYn7BmO2WnUEzNd/ocOM4iUUS6g2vhUhAnmjDXP6MIpGl
fEFlIn9dmEqSfw5FRNipf31qxdD3yOgdQQ3SyG3NrAZ55oxqiiZ4UOg6y9mhSWVU
PPU6L9OHwufrOu7bHJkrGvrcKxou8b2ZQ5G/Qf9EbZPHboubltcGf7ZjgOGzw8SJ
NA67GiKJzNFdYNqGFMHTRfDr1zU3/Id33vRxYpP3FTTzMSqO7BiBOzWiHrn7RWiH
gJ6B18QZFo7ET3XvBORZFKMifwm9xVuHrNA7bA6MGM4xPrxsBbviGs/HSnYgGqXy
HNmsCcD9T/LdC3hlkRq/j2+QlPh2yCKAHcjueL0C1VgNyyhZN2cet+z+mJAq3RWh
lkIYRIXAlKTadcAr0y3OkzbSgW0suKqYq0OcN152ZNcSpDUqISOWlUQohY42mS5B
LWCGZYipgTp4JHxl0I/OMp/tUzJvUldxCaFcjBKvo+Gfa4evG1OZyeafAtJFavy2
AIMXnRZra53iAYP/PSzN6Jc1/npnd1lpxH7JkMV5vDs/HDZh+cfzrXKgdDFozJn/
o+/xTxbNlgpP/93XCPLUkNY9MhaRgp1dOLNNi0JtTQwQJ9uzO7W65RPf4IHI1JI2
Yv1RwQYGhaIYnLrO8orL/bBn8xL8lDftRyHta4JGtKTFhZX0FhTlW3n0NNQg8yQT
FOp8Gps20k2sZFSVNwtdV1IZIB62iyYy/eddO+XPQLU374pCBx9o7pnNHy1brdL3
DDR2fClUy2cROxEz+3klcnmlZt6ExI5kDHpMa5M0u5VZCjiu0irOMWlM0yKBzhpW
efNN7TAduEcG63UTWzN2V+tGRkSeR7Rs8yvubRYpgNKAnAVxp65D35PtN0CetI/9
cnhvACwiJShvLtx2Pysx1ch7XKVk2LNxxZGaiWfAH1IVMCB+OFK1TRoSeiD1lY1t
dANqfNc+SPyairXpTf2qKATyOfaUwUzHsRYXQZclR45xgAAqB8yja2GFo8zFzziY
IMD5xlLeM5Gm+LEnl9VM34KSKw5XXMRwSyiCzM8IS9TMlKaraSWf0jrnAKTvTnz4
YSr4QBrB60sg2UCr2K5CDX6WuOeDRz7m/bJX0S5Hxi6T18VBdCw0rMKzFhNE91uI
RqcGvrU85mA+UQyu46+MnZRXltOHuVVbcZRFZLGxI3A92tJQc0Jsix/dbJEwp6+Y
OmUA4F4gkIgSS6VasSk2Ksn7oXNosZmHjox//VWSlzq53uE7UBxkChtCZpBQyJtD
pg/UM3xMcwpodAbHTUX+H2Pc8qDHmyQog+ILfrXGDyTGDtKT5/7ewD8HHUgMrxp2
qDFQl4mDU8KQFAZGL+QdsWpk1ro+jJurxIC40tCO4YfWuz4Zlk1obdt0fg4EZOJc
wtIUcmq6s0EyZ1B9Dv1vECZxYrmR6bg3AwpeZ1PXdEO4x/I6tJ7gtXix9FMUIJXa
xfEnfy4x/wIWpfnujiCXC7g4Upb+AxDHU2PWAlKbiiP9v0U/fbcDRh/IpXP1D4Wj
D916Xs5LRkM2jzWiQY2wG6jd2y4bESYX7fOY2bB9dRg3rIuNgGfVCl69fXc1xbBT
FkmDEin3a0nyd3+gMNVs3SymqpCPlLO+miL7b3hw0+uss8Ud/LLCPeX4SorhMd4Y
U1YTLtpWBTuD3I7AMEJF21G9TH5+QMb3EiVZTccsP2IuVSmC3RnmCxEFHKHpXvB5
W8I2qi2XRjYvkiGRGgv+/kUV17Rqxi8wszBlwhdr6Ugn6wxnn7YVxq40H4Iv4UYU
gyLFN2bKHpJuQndBHcVHR1agd2iDj/F6mPK/kYMHX0THvg+paHAxm3dSqb70qFB/
17ph4AKd4DIBkdfQ1CVtN+0IW9V9hwbEXTuHo0z+8SlQu56N7Aq1GqMUK6/M8r0j
5go0JZI7AWjBijdmfj8TaRnUlRFnchtFPZnjCtWKNziKStMR97nzR7wH3ruEGY76
VXq3Xg8LfZCaDKlYykxpUKITAAMTW1E3LmZnDMPkau6AKmyJrcA8bHBPWxPpbIqB
DkSOVFZCl8AZAbykutDqYwi6c/mwCTNoORD7HXGuUadRxXG08UFdIyygnY0SqFrh
mNw0knDYssa3td2+ea9l0ccL4HEoFwu9JkonB4yxRvMlE8ybgQF21e+K6op1xmjQ
4ImXvat29irXz5M/LHfZHXvhVtRvY6fePkERVOrRT8UbYpg0mLOP+fwTfU8AW3TQ
mZtHAuZjNKX2IbSAHfQaVM3otvuMFt1AmKhNwIvUVK95YIEJbshWde5bvebjdgiC
ebh+9yw9ixLKc8orkn1jVcmNjN7O0Bdf+onxNjvA6X+Lc4cHSIIHl8NHN0V9mf9j
Rwy/Bxttn+4K+2Xkb0qzyfxpBeTTkYJQgA0pl0cWKD832tF1FQ53+LIZdsBMmRR8
Jr6isfXNq7FnOJn0loLKXerz0Qbhty8/p2JjT8pGEaJthCSl9stTfqU3lUVmldOg
va+n5IPv6Ar7eekyxoYJvbz5fuenGkfj1YMvS88kYGwZ5TIMBsxO3o0tr89mJnmm
1mCCo00E7emitde4g1h5S0EbeTH9WoiW2TCayaujNB/EZ+onfoVWnG7CGumz50SY
ShGGnGZZ2a1NpRsFRzioRMq8sdxkv7SVl6pGB8++Rk5G5t+1+GieNrqgZfqN+hA2
nEw9RhDoP5ZLNTDO5R7GABpZM+6ELbtSe87fZ3RF+cXVYz2KoKVRBg5pLusu+t0R
UElxB0+PN6UWrKy98leW7yAWHz49Bud8YH/aX1ZGFsztAlsiLhi7tJeCugyQnUhP
xCVeZ4vX2GmW5G7ujAiRgSNlNBUnkfr/G1JYQ80MGLsWT5BIcsMRGAt06hei5Pzy
G0ynweus6Viu0Eou36JiF5MNmOrIJHaMLglsnauJ9+PgCpkXOih82zIsp6HfJVxe
A/+oXrogL1bQ/EhfFElG5Lx+lSPVYAVQf/xwAj0oMMvL3f1h1SU9T+9g9pFIy+JF
RoM/THBduDXETnCxKLDR896i8/6K8lEPnpRWwC+Hxya3j3dN0IT2lSL0BeYkj9c5
DfynmXfTfqM1yAjmFJIEfjkW2lRtOPCZ9n8IDgOx4llu7ejNSvjgMmFCfkAa1wPo
UimpNzEKpNH1gmgtDfh7ruEqShh/1iQP4HYGzH0lTAB4f4+lwLFmiRXZ1AVh0o12
+Ock2GlU6w99tok45gY3pQ1d2jkNUURDbNzlYre89xLErKAAO2QVm+RX+BDjbO1A
0myiLBRIVzKJX/BeCHQJ1e69YL8cMFykLl5r9McfpYH2E58evWBZ5XXLC4FvnmVL
0chnPr7uCT6ejDhVNJ5sSCiE53XIp6UPQ5CQRZW66VuulGvtRZfXp5wbAphPXyqn
I/VTCiVj65XIwk/CnAKD7nDcGSGaufcvYiMNaXO4+UuQAWA50zixam0+35ereXlS
3g4OB4PECyIn6n0jz98KWHz5m0cIYLkS6jnaY/4U1zETnXMUbL648gHwFLJFRj2J
ND2UOUDsqHbsSzQwUWoPaJ3A6Zz8vOZD1kEMPavvxco2R5BBNXJ1gVc5Qpbcb6rb
tM/2Rkjv9BvKv1U0TjcPtCgvh01WA7/60+dFVpsHevTSOdxlqV/qz1Z/LmlwnX2r
DvYDXmWF2ooEOHUpTrHfTB8/Hj6jScLOcNcdsEL2S1LX2+yhLeeLyb0fy7tyfp2H
a8NnorOraG8C8xDL4LkPNETBwQKoRMdIhujgINPCM2aCWtGsH4LK9RNLbpx58/fq
IeDqsecYjJB0UiP99QAQGLe1pd4v3KnMWGBrROU1Gl2vlUFEdix3h55BkMmGCblJ
UnjA30KY183YOKl0NStnumyuLIEDY/ns0AFuGpqcDaVPWL62bqhpWpQhVcptc3Si
Q+bk55h4WBSQHdKYRk30AM2FjBMo82AP6pJVVTFcIT5BRWfCFHsvjXnd5lb3OBaf
KDzcNo7n2NL7SEuhQrVk7IE0jMAG9vsMT7HGx4y5CPrnWMLcydxP8a9Stm2Qsrsk
O9/+uqeo6xPrMTrnxOjbOrTVm0vO911S9I3EQ4fnJASe4vIz9oRB25HRuWIvp2c7
qVHsOAX+G1LEYNVgJZDuchwNGOtlpjd1aif9b9k2ATsykNvqSGgFrJHfRMZWTgAh
hfikYzp6VJ95hagptP5wGSolm1CxkbTc1nNyfi/5xyZjt7cYcAH47XDNtxh8c/6D
CxcaMXDLnMzWuNvw5eYGFebt/MCOKFrmc7UKCkUUt6yAfFRZLLmrzdGnp409EImw
jJM5dfzv502yK5dyugUB1PXzI4n4JzLbtJvIKbEa1B9ZCUntt6F/sYitJdN7kqy+
QiwAAkwnIL/WfyosiZEelh4xexMzndKFOARD1ueqUHGXNPvWfSlhHW/UM8966Q+o
Xv6ou7jhyrlrvKFjXkDb8xq9A+SofvGVRZuSmcKz0wbQ5KtcclsITryxwL4lMZC9
me5z07khLudue89tEaJZsCw+8CpNBsHcSoGAkGdTUyiAUq2g9F5akkcSdGEtIarh
rj8HXNdTLC8s8usHRsonNuSuOFr7ZuSgDLZS8iuj3q34nO831ullxiVBgmTOSCoh
zVPjeJQ+5dY12AiJ7VEf+BlDey7eqGkW2yLRTD9lYdJLjAYCfbLP19yaPbQuXEed
mh/ZKiLniRQh1PKFnwywTAqlWTAFUNsJqP79McuPZR/W04EHUNuofqEov87pZXUz
s06W79UCYxPz0vRocqVhFQ3tbxPj4bpmrJNztrE7I94igNFQuo/HK/2mNDkWtOjr
IVJe5kUGkkLmsAdHiKbsks4C7VpK7mkNCEBqkXIL+K0jhknabWxneM7bIZcGiy9P
9DcE/UmaX22I+8CR5W6x/sVw4V/zcYSSCHMKQH9e2xBnEwmNPcstDdlg/LZi8UF7
gTLx2HG5MvG71/GAFJUaBrDq1v3Hu2NQ4IjgZqTyE1S1awM/CpRWrixzLLh78TLv
o8iGBuQaXweNtM+8uZspbmtABvps4LLzlKXA2/xX8/KrZJI5vrIJyqnubGqWi9Ym
51tshpK5Zn+CQ2MWiZ0vohbRXu8ql9ZH7LKrLhEZRQyUoMNcMFw5PFckbxS8Dn8/
9EJFvhyz+kp2OFg0G3lsZMtnTjy6jmUxEA8fEkvgHb7+xo4AINk4lSwP82Hy3unE
B5/VIBmoJ/BURhPGMcOm7ls+EFF+wakVmzjcemmGRFBvlsCIfD0DOiOvaYxwYxGS
fqNctKWjywr2jmvQjj7kYS74z5w4xdQLvFqG2Q1oiaw6PFsYLRWxQg24OLbxHdQv
HGV+OVoB2xA++eNw7HFSuedFxKPkGvD8qyCIvNw+n/aDtLV1tkaK83pc6ufUa1ND
uGudHFdkMB3596MagCmnZstbbNowmF5yrBnL/qK/c+txOpvgoPgy+9A0LYeHdC92
/2LfxgMjo02FVa2bFYwl5jPnhRR8m+Aqu+dBVWrOE200X1fhmKgunV/0xLkozfic
fFvAxkQM6gohw6A+25D3IUfV4piyNUMlrPPMCzuoFGNGvxU+mGp2//N4cWFe/sQ9
uwFcUvS0guM+dzJ5Pv/T16mQKYKT+0vuHvyrqkj2lw2OPyvPXHNt8RoSujiz4zqT
UGhsdcGcGdWTXXYDXVbEkWigJTUfUTXyrg6ZBF/xv0IdlNFjjcaoYx9kXeoV5k9u
ikyqd6NfxhCGBQcfgSxLg0Di9kBk8xYVU01Cmc8/FSkbVWHZAZYthaZ66Atbteui
WsQyl05F1VnM4mO67ZcE5wLPUwKIWgYkTj1C9X0F7EQr9bHYWnM5d0Rrnp+HfFvp
qSUfkoPnU7jlkOyfn0yWf4cyHD7JIIC2W9vwm0HPMczGsHqI7uWiyYV/51afOsiv
dJmD7SLcKF17JgEu6C/Y39a7NYu+AmbHosKRCMgTAWO19lFxHZLOyCWifRcR74Bj
7v9ZochhOP4DxC6keAt7DVVdlPJCxfUhmmycOzz7d1SeiSYb4WDMCZOlNgU414Wa
dUYym2wAq2hec3Aw/kStgxsIOfN/LCGtZa8klhOdTE1oRE4kCSbdNNCWIgoGt02s
GSO4A0rddgQXMlb0Er/joOANDH70MRGrkJEgc6mPTaXPn/nakAFaHt07zJZlF89t
7LANweCqniFgI5vdhlUtv6D1Tm1x2fn52oU/7AorluyX6zWS9tDnznNS/ZYhEYwx
Pvctq6/S0uNBdQNwXf31PcYtgIG+Q/Wvmrw84mW/fo7ObuBwg2wXPa0mXw1OGM8r
WK/LKbeRVi4GGWhAtVr4ojN0sQAK/+anPAsVVvv7pd1yaaN0MYfGa1Or/YBtg+F0
Iw7uO9anogWSbaRVpgUDvGaHSDXyIGcPblrjWaMRFd4v0Id6YGWtab0wrkGHnNB2
WqPXr8tY7xqxy5tX8smlZhdPrNY/HvG/R/g0pHVb5Nmz0WZA7ecpkQ/4RLd/kKtd
evEYQs0zSvlSTEGlE4MaCktU5MRbLu1PfMmPwLs8p+iXsaEOS32tn/6JfE/NHxpO
M1du9XMqbLgWaHQX3RdjOTBBUQwndYWcBQQNerxbmfmdeKlSYxZVLzCo531WGLJS
PzdCZU3OLblW6mhL9VEerQPcRHqGEyw5VypKOofWXXyxEJh2thzEeIZEOIWE/PTG
YymHpbySrv/i47GmUcjzQ4TrFjTyVNbKgaVsA5kSKhz8Ox5vJrvBOKD4qIA4hz/J
7jg5sr6gN+yM0fvHMw2AabQAshA6Dwl8XexNRaQ/xjixO3M03/YHSS+i2ojehMmL
TYJdDqD50aLaUdJtKfOqFhAtlEsUquPIkDOh61PM2IhGwE5diEulKY7/hzrJRhvZ
V0CzMcN2sTRh09VIB09P0z9LONc/fSig2EOSah/EkBTP5ifgJAi8DEZauh4V43x3
3W1CgWPsIJaR29iRhthVX/JTPUbG4sopBbxxywxdDFd4yWBrCoDf/MBP357EDYm0
4F2d1P4MkE9ZwOETDIV9W1VncZEdVexAaHRmOIaZ8rZeBACxYfPl7XrIHVr+S451
Xa5LELmWPRrD8cehUQuB95oawIIge6R4mlZp3EX84TrqHVvNp8BWWR3fIHyR1G4j
xmXTORsz+H0d2UMhMFkXBC5fxkfLVK/quysFHmXZobtkPIHpcEHLnPgMZ4SuroKq
74ORofKK9EsxhwXqsujfKc0tjCmHRH24q+omEJ8CI+SP58MSoYkmG9tYSDN38oyq
otwIlH9rkWvq5KdNgaUUBXjnuEPHEvSqPiyN8n0esGbysE0+8aVSaW+81seil0wK
/F1s/y76uuJGHOR/K0Xaq20fBXYrwhXQOq3yiL2ZWUFcNw32WzJAdTe9aSbShnqh
+GOUA7eWmtfhyC0MVj8XvtGjSFgZHdDTCrRPTCY01wtMwR5cXjow4/pmi6HkcdlG
MCqUl+Vu8LYGPgQ7zHtZaThkPGqIgZeaADSp8fvkyICFLIO70liHyEqUnQdBSgFu
7uXi4vQyDdHS+5tqZZbCfa6ZhTgDjXdkNwMj+puyEmHkuf8z9dlCBE6sq98oFXTm
Qt8Ysbe4RO4/OtnxEktOCWiQxXxG/4keJcdFjAO54kmjsilLlgxnIuxa3Ec7sXUz
QOOkZs87X1v6WvAL/XnGD0QM8DtBQCdpHth23RCqdYoe4w76FKufbBdg+8UbdNxJ
mF/tj3C7lM8wrYrAjXVXp8HL7+AmVt8Wey9Qax5HXmlK9+Tid2L+i8AZSKlQPfjw
l8D1rwhKZmZ0Qa0DFpRKndRQmRP1LZ0M7XcLMp+SejiqK0qLRQ+pziK6k/gBGf9q
F5nvrUAhkO6SdjQE7dN5q/lS0VuUhErU4oqFeWSziA/thTIn7X5oIfdRfyKNDj3+
z75ys1eg1XzJ0xgfha+i09WXwiu2uzL70Z2b1Z/iwlWPt30AePcje4zFQomDdQ+L
wNM/BdlY9irSsdujmdr4CrWxeV2BdqswfDOWP558O/GvmJna9u9GySi2Q/NhX9FN
zhVlHjiKV0grTg6ZNh7QqGmw4qxBu/sfe9cxh3lvmV1MZFyDfSHS4N2G7TzxyXIH
BBNqAlf1iTHrk8ns8uTbldBumJYjr6qxKxlSS3UExdgcaZ8WW4+exTYc2yoUK/l8
1Cb8arhKxPuposwhob7yciUXruawVlTQVubAO3Gp/zCxGqYmoan1HMnAYfb0HLSU
vLB0bCiuzj0rJKCpv7jx5bdshFgmKpVUELyWlcvE3fXs+D2wfVI1Cg24+J9eSCcg
fEPE8OPNpAaCBJXEqgIQ9yuyMZS4w1wqSHVY5Zu67+W7eKkrZ9Pr0y/IslxIumom
vvQJIEqxlIw08F/R/E2eFeNFcy2yYAMvLdGq/IM8/wiV91wOWzJqRtbWmU5cJ6eX
QdO7+Ur5rHiEdXaOUvChVF3mbMl2vOjQftDaFJp6we5OcamsN6Rv9Y2j3kZJZxJV
3fvLlyUV1UWiSw8gnuU0XPv1WfI2mk1oqvJPgxq8PBNGcuClUxAjIfHq6xvEHOmQ
CXWWFJ3VMASIh6KBlTyyUyweIr0gbX8OKwRuvVq40mJ6NRDZwmd04zEYFw+qcwb4
bl0AxiuNg1gN9oJo3Eo969+6t122qOVk//77zpMxiaFZDGzxVuzfu7wJhJk6V4Ci
e9MhoJiuZakzkHLbnOlkzaQtlj28NZScSFP+M00b4Zm0Z7BlhpHH5uE3an3Fdxkv
qPln6fu22BnULTmdoH1UyQs3RkthaVlI0Qbe7CMcBfmu/ckJ+jrkEg1pDrfhJ6jN
9GSPYOIMhS1LpOywSI7rT4NeG6iVj9ZcoNNTeLTSyhQ2q293CCrtVeNjeZbnzKLs
i2WsxxS+t+02axa/F/5xjrgHP18L5IUegjfoGitIITVqMoz/p3IRpIwnWZ6GGl2Y
Y1rRd3Nz+Otb5WcOq5k6qVR8aKVB+XT2QhHiTodIJ2HI7h0YhCFiWfO1XX4ydjVt
0I+aRekMuK4aT+0ABQfPJ7eXUFbM1Uvn/nc1BzzbumzRxUUf4wERwfk/uHxpwTkU
SmgCc+hCC8mkBPCwhqoPzJRYkvMZE6/wc5EKs7bNcNAIHGv1pC/lvxKPGlS1wsde
P9fwWXHermdLVP2dWj7b3eqsOL6hI67/RBAZ+fp7dZ20Cam0KKDIS8Sz0GJvj5Y2
WhHVrAfQpf3N+vmlqpYrIN3ilZmQwiJDjU3bKySNc9dUIc8RtklVZS9eGgvzgISL
DyWIeJf5NtGDB+NNShdb3FmE5eeBnWiAsvG+W+6IcMU37ov/mz/+FzfDa9ruFXST
hQGyoVDtWsGOuTVa2/cY9+NWjvOKwpvG1OfEbL1sX+56EhUC7MiTsdq2Tr+boTMJ
9Zb/gcx+s/1tyrnqqLB1EckZLlXQ2ZsxBC/jyChKCXLtTgSiNyIQjd4fLMLAPZCC
cQkupTsq45QJRf3tYW4N1AsSU1xzDmolsLeuUy/sj5EeIzVygYYEkP6agbn6zn0A
3hG8z6xaII8FuaSLO/Hag2aRdjKEcNPHPoE13vVIHF6z3SC/oNlfhxI9iPzny/wX
1IXUgnBLwcREC763K6TwYnr8s7S7v1CNEMuFkrW+Jmie8E6VQp9eZkv91fi2TkHB
6C4/HipfJeG3f60UhLnTVfSF+GN6ICYyak3s4WeIGlgft8GJGHiIRJ0t22Wv/3Do
gQAs5RLSafcaf5g8zg80WEmxBDJLi1v9O9TnFmswY6HBaWYpiRcyj3wWuZ3QJs0Y
J1dpqsAj13Bc+YYAchNZCMZp941ZnxNSI6UufTa1paaTVdmwuDx+HGjDk/PFXDvd
9w19b4f0eG97/SbMAL6GJz5g7StvPqvJ9Gqc2lw+5FPMTxGSeMVkMCA2wR6kqWXs
Lv058iexfJpwH/4cQsKrrY61skXnU6OHGxBX1ijdAvc1/c8MEojQ0SRGpARhbyqp
EL2ek6id7MCYUfYW+CVHpAvhH5svH+kFz/STnVoAndL6+OvPqdnlWJ/AZWWv/ya6
HhAHMLwcn5xCLx7IdPy4+HQDRcdJKD2RIXiS4CSX/epLPBvfvgDEVii/Oz118uWP
55f4DRCm9h/x53V5eHZ6Fuuj7q0oMBffDcdrW09LFlabvpUAnPhGdEUpYZUoctMX
SDthmRV3KUG9k4Go8FZXjmNnNJRcqEQKiySqzP7QyXjQkcIpbMJD2YEEygVrZzHx
xPgABmSTlkm74a63pJn47cH7ACuTREkENyxwsVj2nkc1l8jipzXc4GbDnAXsD2Yp
pU02LQsQ34kPXZ4GyyEMajT/CIvee3M0bAHYA+irevvWU1yUoy50Tgegb35jKqoz
dP8/YNm2RhddheObbWGMztD1kUMiB3QCTk22aiCdlaexPaPljUpsOVkH77vZl8UC
ahsEXXzfGMddQRWMbjUcSby5zMn6GifxiwOtjdim4/cA0b+d7etajHBoqU5TLAAZ
ENanRTQnEzn7wnVLd9eqNBD2TAgqGdO1kQ3VKP3pMnmQEdfH+whLCQ+aYeu/RJg2
NJCYQGl7emSjvZpxvL5ynoS17+aG1RKVi2eAK6KP+l3AaP+R3XjPfmzM+MSUFqCI
oai3+De7qX4dWzrTDudRFjevlh0z1OpbHIqGCA9R4JgLb66Aso9nV6/AZ/bSeR15
mrxeEu5mDxzKuCSHh3SUAMFc7Nb5X5IzkYoHcSTz56i4+Pg5wwlWNIqx3RAejlUm
ThcbHNfwT1ySOd2yvIFrzswnmyoub/v88Rr66uwNInlA7omqdAjAgnE36OBsB8/7
H2PsNl843wbn2nIfUvJADaTJVS2F8gl6z2j9nm2Ia/fS682jgj81wfFyqme52Tj1
eu8kt/0VLf8A9q2CvhGlPZW6cbZhwCpQ4kOJnSHcWBVTf9rNcSi1MB2+02j+vTIt
Sb+j36ItMEHkIuN/ddzp/OhaFFP297pQNC9aA8M1x1sZPVl5E/uLm/7ExoTPjG/1
gcfDFR/phOfOymDdc9Y/2M7UU7V1XFwfyEfe+AK3oe7frnCDuMaOmnwKXJLEM87f
fLzu/TlNP3ImntbgLwi4GzUYf8oLObEjhTKklpMHs8+2P7ZBHzP2ebVsH36qztnC
4UzQstGibxBLcxV6ZneOj4YtI6VDV8mN5g6UQdqieXloXg5idiuo0MFKSZIMt4Sw
/mMTRaTnltXRLJZT/Pb69S+sIZvwA3buQ60J7+fEWMT9MPXPJ+3G5JkjAKMkeCoD
+bYstpVbFaHUBaXSsxiZmcXV1FY2ySJKPQgrufa7YCgxPwn59kzLN+8UDhz6GUdb
M2/WY2TuDhxFJbpPkX2BUfOgsrUnDjE1cGgsnP/rZX0a17HHZwlYwbDNuVSGknFU
TLOqndaNSvbdLqb+uaptDCIgjXk+lBLdXY2AD9ozI+VutSo/TaTtZJRgNELxle2P
TV9OrLXUSryHpX/tcViAnm3/wLAvrZgT7e8zLFNiSvHLmwSR8JZ3GAIH+0giduOb
Jha7I7mxaH0E9i1znFh65AfoHNwo4dKXXISNtUNbeFoUv1nS571SEoXDiHBRUkHl
rwg5XAGmt20jJH24PW1HIXat8ZhkJ7+vNFKq1c8EJM2wduWxnmyesWs8nCV6tcsV
Il79PW3Vhb1cOFzckxN331TFJGtnUH+DP9kWy54zAl2jbrsHQMTpRvcCoPrxjNmk
UMULH0eKASxA0Oxo2+fC9erUCRyj92SjXeDrJB2U5o23puJd3X+/4soVnpvbiPTN
PUN7yXCQAnMwo/zX7XOsTlHyd8ppL/5ceH+CoAVbPqduaQ2xxpu6ipJjWwHEnhkf
ZUU+vLoLpw7TxwwNifbOfamDXWZ6UAG+2I+T4z2WPPkhrxTQJhgEHVRI1kKXccOp
UGFABrNgLh1ai6BZ66bJgKrXMlrXkcU5/5p0ji7DeHQqwsEahQ1EeOcT3Xo4jI0T
aDAwAHUOFDutjY1bUE8/K/+CodUANu3ArSpe/6GH8vjrgvPx89F/CBdsfM0WQ+1S
RqGIXdpVLUtONL7uySxuI/9gpKukYFIgUHGSOse9VKv/9fM5a6XWTo3BsQpJ5Sad
HdzM0CMuDuDUikhd5HI8t34UZsYUTIujd6WWAh23GomdNqsZLYNrU/EBIJl0ziex
U0NalvIV6vKU1Akk7kqnjWIgTTbPYnKZTpY/wswhfIQyi8uyNs+vfeDo09n3ETyz
6u8nvC1agd3bk29+cq6DV0T3/jBUSDhj6H0j5Py9d1s+vcOekWf8DUSXgIdFRNvC
LJ9dMafz5nK0F/KTevM+TetpGT/RzBFUAdplwRbPjLzO0mj+LAHp/pbqLafIB3KD
jEum8wP5EsLS2fi+4yveHkxPq/Zb2n1ajMMmimj7CvgPqTOaMsVcW+eiXHvV2kLS
39/uJH3HM3uQYt60uEHmyEpW/GvcmDuCRQ/Ve0kRQuMEJMxNe+xl2ALZzJx81RU2
LEvpQI3ZeguoFQ1kGbwaRFQXKoK4vDp+39wUbXo/UUb8MuM/smPZo4AzBrUGm9Fo
9yMTaBoKO4SA0AvEYxp5dCP4dFf+WTqPkhPaYzlGErkHMAcSCk4RMhniW9PJPL0X
+m9FhlNGcsy32itpj8A+Gm+iKCmiQdUb4imiCbuhu+rwZDqZVmBqwn0m57akdCfN
aNGKCNJbs3ViIN+JKqDs3AgBW/VD+7mB2FbGupqeqNJLtzFM4jS9Yb+2p14+rW3L
fjdHYE0tNycvL/EGTsEy2ag1WLuBcn4Ndl+wq1ArW5OabPGY1ztM8ORUIzqkHlwq
LZjwC9jOsj0ml+90XsJtTzoDuUxdY5+eyb0LCqN5KWqGMvnNkro+i/5molDFO2JB
N943NyBQJVfSUqTId4HfknfIXpbW4N1Pl7b929IwhV9KVD9XMskPsm/Ey1bOIDwp
59Mmhuz3AC9/qxKYfEVZe/D5eI0D/MpwfFrvpWkWAvetdIOSARFt4WH2XsawfYuz
apYpfvKhGeyzS+sur7dE74oIGGKffTRw8y/G0vUd0+wGsQuRsd4bWwfGibTk3djg
7rAKc+DoC/zv4VFhtXO4uFiAQoEdI4TPH8U7+5FrjKS2MPb+DYKFzcUz0t0EeaW/
SMiCJBDqMisGfMXhEyiWu8OwOLl+BuyOdEes5A/8eDw2F1Xberg8nYmRebCYlSk9
dSnBwgz1rip0FFkzBEQ22bN8in8PYw86rUIdKvViFsr/PV2NjHbcqB28IiMrdIZU
0Rdq9Qz+mIc+4TEif2XHYc3fYePCMwOzDqwZL410nnJVQqdCzWR3Vxau7fc57/pC
BTNMNnJWiW4EWA3rdqg53wSJyqxecPuj9DH3wl3g4QDkNNu0kUIY+3tJwMMeCVK5
IZ5/n5Nl/fJViv+R2wWssqzouN1xA6GXBaIMZmZAtPVmCl1OowTKazuRCHmV1U9s
O4guUCjmtcqH2IbHBgId73ryBs1jKxaSn39GhGGdKtEVxy88Pj/gSQgtcuprmy4r
/wPN+DqzGcGe7y4vrbAal2bpSvMGUOueopGjM2MEJ2RNadoqU+D8iwjEvyLbjPXv
2riVqZD8eQr+FoZZfu+dLvmYSIPhuFS2fnyMIsgEXgisCSAvAKWQuqZlw/lbhiJ0
aanLZVcmi1fJ+ZMJR+2TUC6g8nQZ8rQjLDCQDE3CFHPM1tcaQZ6Z3LVv1ujnRX07
vLoBq9i0ozQZ3EhcfupYLSb/HwYouKLQIDLI/yZDn+pdRpi1sqTxnzTSukswn5N5
CBNlEgHFH5S63ni3Im37a6YJzoyJqrTvDE+hW1E9NcKPsxH6V/1wBvqBtWqt7Gr1
3fH1ttXN5Ub/oRP3b/+juYQDZz/OeKNTD8jCVfvRBGknCtAA4AHJzcAYER9EM+yr
K4T6MR1H8yn95ryVLIdLUE5q2zRpHu+23gKzX3IhD6zyxPIQ+FcHLg3BH89Z9EtF
W1dgeNkrw+B5cYHDHBg5S643pQ+UArFNTb6a+ultINmDziNPoBFnVAKiCTdA7T75
GfW3QQEWtB5z7TlvilEbsl6mk9HWzlMhhLaBmsjLC4fO2VierAjUv8uVSKpuH6CR
MJKboUoTz5Q0Oo/u6A9GBsa3uesmFFjynydzNz/D7t2aksXpngLE1M/hsM3zPgNS
/zj7Y7mC919u2aZfNHyrX1WnE5VlgOQv3WrHYLe20SnF2zX3sNaGVhtLbIGmmJTC
AGAtBTs2924OOcnxLKW7MuemoWRPJIe9nvx3ctvuNrXRpjGm4ObIVtUur1Swirx8
zYxD8cqyBxwGNFTTJ86eI1od5oO8W6qlEUoB/bJmGZGDEz0aQyDSqhV1KJI6LRtZ
/+cmIwVnAURFOQf7bbKDunGKSyvjnmQNqUvrRhefESIVF8a2NGZMQqLjhcrWkuIT
DNnMG/TfbCHnwnuwFiUnset9Fm/4e7+W0crOOy0QpW2WMMDM+GdSfyyGBb5r1ydC
i/mR8JvXmcVKARogGjKOLjMzAN5off4yqhoCPUmvus4V/bGiC8lmtLjTBDZ9c6mq
DelEcucZoOqnU792D0WT0WY8BoR9EH3T4WLmPe4liqPkWMHZ1ZeeQmKrOSeHPsAb
BGe8OZFSpa6huTgW9hnGxH2Z2Pf0Juofsbcfx3bWHnfhx+FXvHsAjVoT8lH0ACuG
oUFeHJBRlDvj3940iYuTlJdKgYcIFkBscYgC2ZNWMtna8zZeooSs3uHIHmV1pLHA
XYPBAHML4/jUBiQ0qzAxHwjbhy+30F7Ti4qkg1f7T4MOnCM2UEfjEQrwhNTtt/wY
WcG3okCBsYmzHBJYnv3PjRxrYFP0Efyx7mMQv8s4UD44BmUjaDarTMnQROScYWoI
Tr0YAnxLwM80VKbDp8pCC71FTDjUd9h+Vo/ZZQ0QowGGoLjavxSypK238pHr5fvU
NTO3ZV81asY6iMb5EpQ3PTLiH/StuFQygnV2DLNCbeGpTV/6PiOu4aytIM0e8ieh
lMaWjPd3E0lXizizyd1GdAvGICy3ZvHp3UrfIBsD9L5mHh7fKrZLloOrmHo7bupE
K2Kl05vAWHo7cILQUvhlKJATM07kgtIjEF7hL7fHgBGlVXQgzF+ksSdOutv025gw
bkMASl//rBdi2sJEQ7uMYf1lpfgXaBUibIJiMNzOYx6Y3HXDb8y9Phjb310F1ztu
8T9lfIPPnd7cnHz9F+0hzaW8c6OsU1aELvwlZdOXOwW8fV2A4GMdSM7P1iFcsNPf
wQc2Kj4JYH9EgF+GDa0QTRipcx4mhNFAlmzleDq/A9uGDzI5jT4TR0VrFBVxH+h8
4hhewzsYhxPtkmF8ChBlz+p7vAhSv/MrWenKTw+ntL5dp99v/TTMR80vsfpPcfUw
PQ044BwTwNbZVp3cZhEOFQgF51yggrKYto7Njj04ke0gnSVwGVXr4yHh9rf5fwIk
fXSgQ7Ap/zcsXxnTax1tskvTRO+W8vSfPpzYfxMCNaKTldhiI2fjExVpz7wqXSlg
YJCYwZ8QHBcL4Hr/XGPZduofQNxA1l+lZ8MdqoVPO6fyfBVe/Oi8UELpkxijbrF8
caNg2toTp29ey+Gtc8BfT7xXdWFN40CpDxiif2d41Sl5Mc3o3nKETGVwqMiURPOk
e0UJ/j6LL2p6hgfHoFwY5wwm5Za0u09fJO/Kwun9yEj9fz6ioYj+aIyP5/BTnlNC
4rWuQY1LOpekbqUIHLlqUKCbQ8RvkkqkTaaTPHMZdiZHezOYOYkoINaOhCqKrHiA
YDKDxtCBUu72czVbOUXzfzhFhZQopneBqcIeQtatrRIBqhvASGy/F3cmatlhxEu4
fXP1UJgsg3yvqups62vB/C8I/YYbSKjrg3rv2ZCl2yx0kDmJA3B0Sz7wCkYzQZfo
WyfF7tTkbLdRdbPyxZpMOYKEZR8sAr9Vr6/ObBt5RGxv1vO6CwhtN9Wt6id9VMHF
1gNXTqcRI2G2ajDX7q8zlxiphgnCwEq14an9EJ4Es+4x/vEOK34mf2PdC0ShWAOq
ReczRp1OagbgaZsHN+6OqkdAv0HXQy6rrRbkdLowwadFHN4ijNykk7unhTrYTujh
zex7Um1Al30I0ohpLtjWZCnKZpGM5pZAgQmnCbyVCoKJwDHvVc4jCRfNKF4NoiiZ
pEu5jiRTQz6Nbf4NKy6Eu0mdG6kH2MDd0Q0nA9aQK1Ys8js0RykJ9k/v0paNtRsD
P2T6gKUxBa7iM90VlN6xhOhNRgFLhqW3gjnxEe5LujukSWaH9TuUk/nikHABM+4N
056ZXB3am6x5D6PuoeY1OX61HFyHAaWyd8liv1nmkVs5QWQO60wCiis/uT+76Nc9
xEoPyTI8gl0HQFv4H/52mBBm5POfV9YyjZYU8OkHU/EpuAGciUouLhfiQ5PZEn1n
b19htXpUHS+9wcivjEQDNpRj+FafhVlfPzNS53JpWR+GeMVKcGQLfFACSqqF5UaZ
nH7e4J3R9ajdImMd8LADl8vh978+GmXqZwLdyS8wdqyqkKpnUpvFDaKzuLwPHvCv
YchvbFy6L1IdrxLfbjKCy13mfYkGKjVlnkO9tFbjSt7lY4MYcht0bH6ihVvVwGjR
pLkLSM5IynFKBW+WSyPOG9GBqBrYIy2fOpugWRC7qxUWSJIo+eM1NIDmtk3yJD3z
SH2HV3qEeT3Vx2+0HMD7hHig9J9VnrGqdvMtfM5n12+McJYBT4ZntK322V1sb3t9
abz/2Gn3xSW0gxsTGuOfE/iL6L0XSBqBXgFyeYeuwJwabC5q2X9Y5YrX4pZAM+Ix
fcqYdUvj9aUaUlDS1PWuw9Ldf6YTIWqOpWHm0tWUI8b8b12eZxhMJnBbi5HunVQC
6oyal8cItIfIPoLuOe5+vjo846YS5GVh8Vs+uGZjplO45x0VNqoeIl32uLobUmCw
QJZtU6yhHZqZnD5JqrbFYsZ2ywt7fi5Wf6gZIKwNFf1WqDYVqG4fYMlev+aNI4HW
99Dru7UU5x95i8+wgXVjIVoiDgdK1G6PJvx9TnvmuCNKgHdn5pMPsYPawywJpYft
m9T66ERe5ru6Xig7bEiMd2uEfZyxryowbMOPERbmIXrMAze8NaPp9rBX4uxCG+XV
VVz+CPYY/3BXjCz3jgp4GXqMybjfBptwZzFKeaid6lKH7doQ0Xb2t/W1/OHmZtxh
67w4z/FGaloSvbsrkRJ1Lfx0p2mjAwdCQG4NjrZ7tiCeCDAtwuvB3JqKUBX7Ac6C
TxWv5LyzxaKIV3fjZ2NjF+PakeAtc3eA2yDQvoFDi34jYYq75OTmyE+yoQko/lvO
kWlB/QsBOM3wXmQN9ZC2ERv3DanfZVdgi+xJ+ReknvCBJq22YEtJbbmnV4wKr+LH
dUx2hCMSeqsWBuyg/9QIakoIflZ6cskTgVt+lw4vIopvBqPRgEtJk43jzNl2BRTR
Y3nMvxfWwBF2aTGb9EB5Rj24w5KDxZpNItzgUH3OEEzHf2iQRTImi01fnVkthq84
Y0ZiqzdYRkvrmm1xVH2EZgxQN3d5EWSunfQIDu+A4gLG8YeFxr61+IICTa1N2pAT
J3DcARmj0EelzI48xSKL465n0noZSxzYa87FhvRpri8+ujJRc9F6aXkN7wZ2SBXd
ZyWHVX5FoThfVKmll15AtAwRBnRRgP5y2witzeXgh0uejoAXrzpahr486Iw2ziZb
B0LAy1J7b0S0ph+tj9LXjyzaSS8JbIx26N0gmgWZsOhPyKvXhfd2bWF0S9zteXMb
aeDtlu7AjHVWlx23Sm8QaNfwdZegKwgJHNmFwUDQmslBA5x5rugeb75sD9A+Y0cz
T5DzcbKnB5jkTRViKCsM+IRpG+HrlPizo3VH2yOAsOCMS6RYjG20Bn8y9+foVQzn
aylQZsIPE5CmAn9nyuj/fhp8sbqUNgwmYxHaO+JPaL0mlD+IvQZB51BMkU0CSvvd
+fgFFSRxsU0GWoIJNyDp3WnUqFp1jPWT0NfjIAEOwc+GFz4WTBG7lCzrVA728lU/
0sEhamP84VNNRf0MQ8lVG9P7tF8cp29ALfm/wsvMgaQ6sMOgJ99DKXnH+opuw1/M
+KNrVfw+Jh83YIs3lbRWRDbg6rw2w9mG27JNUeB3eK8NVlj/S332g3vrT8JyRNpN
mfTPO8ARAntu4kfyWHCZTqcbJ0sTw8T3nzrTKv2FbR3F3xz7mguept8qqo16eBkM
tAn1g7AxP40PZdXC1zbyA7UiOFgYGJW48CJub5iVtxXRRxk03L12i0mFLrqhV9pz
9cdt+KlB/weF9xQ4rM6WZCZqB451CoIlOII/HizisSka0fdT/1xb5tJMbzMSJopK
/6FaBFITACuAv5Zgb1KythRlzmgBHj9nQPFehbOQtYGeHWD2yEFDwpLku83EKlpZ
d2bpgaD1duR25HO+0+AWoG07mnyjJh+ClG5286W+uTcjiLog3S2r7xJCdDUMnPGP
KF2leFSaEgIMjMwPvZ2Cd1S2BNY1Ub6gkxM1/qeZXxZnA7G7iEgvmoU2WTacZS5W
N/FAYaiZpIc0WOuJQPXn2XQRP3eTnRRXiKE6HGqvfoNPXO/l97z7rTIRRW8bPQfD
GsT/ZgSoMN/4IiUBb3rVHgn1KuDq5yovvLCCXOiY8CBfQkbiF7a1iCjEyMHYT3WI
ewxNH4qmUpyth/YiARC7USRb6/epYLo3hHueZNDZsMIy+ixgmqF3GgAHKr5T9gQ/
/nszc4kQm64CdFmqnbnDDJOVjB8yPJWqyf+tDveLQHRmMCV6GIAeGBoSlaAPAJSV
Uw91AmDD2DRt2XaGcICBDucmWTBRaRk5bVsUVAVLrFPDHI46hP56NmynU4lkm3HD
nOpPoHI+vea0mjkh/6SoyPN9/pPNquVCzaycjeGRVOJhEgxf4NiUCN21R2bTrAnW
f9DYUcc8UrnQnatXong5XO5cIt9yAh9KecQL/SXIeRkiCdIkyYk16J+wos3wEc0/
19GDBfKibJjnddDN3cYIehNk1TBzl/VIM9c/DumVN+AkeNC09wnv6F12UMcQGqrp
vsO4u3KLZfRGT5scMICn9jZr+E7DbzCoWuurSFm7yxGkcmaqmvohvWhbgE76jZxi
oVQXT13YdeAydwDK/9MQnWPhDjoqpk9wrgPPdxOzuT/dZduhPhHC5EACyTCfV80F
+rZG39zNn2PRoujCDaWza/937jQ4IOCo6y729u8dW7Nhzxw2KTwYg4pifgvZYVLB
E3g1lHgggx9qF8rzFJIwoCFPMHjVNyX4i30QiLY784gZbBTwvuPxC48C1VEVFrbz
rllF5F0u/iYtb5nF9wIM15erYlm+zHc61ioD3MPuCepfrJ8tCjyAdYHZC3TkcUsu
6q1P21cDihQRlPSzg+kGwmTF+DI/dflp4E72GM9pvHpjkGna8ymstzxvk23Rf/Pt
HqR6/9U3EgO4NT8G6niKUwKFnMPY1aiu0P/x+JdE+jYv+okjWTO1GpYUdkUcWcfS
G4ry15RUi+c4dhwCgPofxam3UeqF121Ll2un1IIO4SShAkZhNSoFO1gkZlgE2fBK
QObZADVWVT5ogUd9qfVyqsMy39y593e8dlucu4ETCpwmJwwtl462Xl31vPCxoc/w
E9+PgKVVK+oALqULRK1rAVE4fPagnl8p32Sfu8EIGDTgb2Pd+F3bjHQ955G8I5oz
Yb48p96EI7rb5QML8HE4mHk2WEz+8pKTSYRRZ5iFA+d5HLZ4Id4ehOyKm0T2Lc0x
QIrTPTaKUb5swLU+udjVTx1uTdbpxHVoxC1/EpiuqvP4cdDEOICIDG9TNWNZpMyl
l5cieWSQzf12LNLOpTtCd6gEqncnbpbOfev1n+wRj+s8yKczCSNHB6xKIX+CGZ9Q
tengT1iW5JyF5z8sXXe+IlI9T0yoacasCNp7gSHws98GV5hh8LsVs9IgdRytbD/E
96JqgYhNXBnO9oI/X2ZK/rkFSqvexrma1I+VtATyBPYjYn/Jb7S6atz7sJXd/wAd
TUrt6MteJ6osSy7Onptjb+IxU3lZb6TCBBEqsiNg7oeTDbSr8y9xAO7NfNkmtrBv
3ayIe+y9hNcUP3z/cmzZPLC6ESGNk0y6lZjjr/7snEuVtoD7g4KRTyDZDVXmDHH2
TdsYnbwFMWCLwkNGPQK1SNvCeicu7zFSaZdwdw0oGdQ3G9q+cYgUbO/PkJWMZX5F
KTutymw9FR6Zik81oVpvFs4AGvA2KQ755dCe2ePKAhM/yXJbSgqcEO7FATlFv/oO
us1GosCRot086/kUy2N1xO/A+fn9qCWmn1ga+MDlW2/wZeH+6XODVl+3Bgsiz1J5
1uYgJk494sRHJn7GQWCQC2EKJGK0q5LU0ald0lHbdvODwbUeLJnM50hGoLrW1iRB
iPciWsiUPbYscW1ZLrAgCQuiqGI4b6gMq58ZkvVMKbB+eqbXgTjTSF3HZzTXU9Gp
PyOgLUZSbUoTRP53NS0SjKv31tDmSPlO+7qJYJg5X/VEMQa9KM02fp1jBVDhyv33
o8/HVYtDCsM3PBfCiYHA124TTgfyjcG6vD8k/gie6Gs48asmdrBs/lunYVmC3iKS
CevOqd6yMRf0l+0RreXitncsjqkGWeKUbvp41WLRPkb5Sbr7J4zazf+h2WLIbG3q
wtUvxuwqr+KUf6skRhwMWbBEhedIJ6vK54udaIpZsyoUZ5r7s7NfzM4xttQmeuWK
Ge8hOr4ZjlgcafDhIzp68iWl/Es3mVr8pHLbuPLEl5Ru/h3CZFcctpUXYyujfKMC
wEOF+UlOSzDShrtjb7eOCoHLsNfu9pIsLCy7qIozsgIP8jqO1uWym/qfgCUjkKp1
PDBiddAEMQN2taBgp0ZhqpUE53cnqyvmQ/UoM9aoKRrpW2NbNB8xMvfyC3yvhiBj
Rrn8rgNnuN71cB79FQYZ/R8QFpL73OGnBXJ4slUXriqT3yCUbC2o3Gtx9LgvtkWJ
k5FuFSbu1HxxPOXyfbZhMF6HL32yDDl9B80nAUVafRMp/Odb1el3yNaFT08/exp2
bFV6z23HbyAib/DAyaSdZGka0Fh0FC9aQTbQ+WUjD7MbQa/tJK8vqQjk5FrORAXY
e/FHsPXZaB65sJ/KIUZHmM0uDm0rc2Ic8LT9/ZI1JfLQTTkM483LC027d+KgoAuN
5I8vNU8d1TJ0gneS/2eIAaq2AQSqU+glIz5GVsQBJ1KqfYLzXwkUTip79IiHY6oc
u641GZczuzGKro4vc1b4IiQtyRzzqigqHYwFuY27vuRgzUT4h1+II2VMQ9Ikjbyp
OJcXU/dubXN7QNxsXNbNjpGsJYvlGMVSp/mUOLKeN+x/6IFL//iLmB5SjX1TBzPo
vsbdvpTCJwSlyemjqMJAUVZNwbM9LOralAR2Rqjpr3Qe1Gk0vOzZGowuxGFZTXAP
jQFIACtvOiWmisftLxl4bhLy+mVYDlAEfnOixuGlQOpFHDHWS4XIpjKf8K+DQMNS
ABHEGsQ22HKfjvLo+4LKfDnqVDH+dAPKpFT79ZZ/60AnFcrh6EC1New8hqoFxxBJ
lLtzCQ12vdbBQHishGyWB894GFD4DcjHbDwHmqvMjFaHjcj2+Jz0NahSOsV2bXG2
yQixaHemp5pvti/0pIVPKfcQ49GiabEQ08R1gAMiuiwIPF/GusYreqNAiHC67DIG
zovcy5oxqBqt0YpHUVs3tDBEoFv3pq6LtKt0rUVEatbQ1ZIfhdLFbbow+UZKamr9
mKgRxlgbeFPczAMukBMx7kM60tgdnsqWTvV6sX50Lw+4Xv1Hozmt0dnENkW121DL
3W02EormLtev59SsgygWDis/JyMbgoXlf6+gEheAvLiBXltBsIleiVG5qfod3MXt
S0iMnlnJopfEJHMRS4P+X2u4wXpuhPo/9Xkis35vqOtIjCeQV4rud8el6JenTEB1
/8uImbWLGWa95etImkOdw1OyakxNkGKpM/mQBAcRauvKiGrc3P0Da9rHHmHMQs6L
pz7eT32R7O9JFhAynn7FuGO63lv9RCwuwwVgLLUDgz9AavzQTVcRTbxewhwJNiGR
7dEvc7nO+CslTScPrygQUCVFTbii5bT2SSq+xkUV/1ERaXkM/vetDQD6362nX9PF
IK9G63vGVIhH0OXccmA1FBWRff21BDWJ+NSRTQquQJoZLaignG2pze/a2ygjjimI
dfZmrO4FdohN9BoQR29jwXfrORYOTqEmA3gcL3WozCu0V6dablKlFAq6FcKDtJFJ
4XEd74NmAdfI2bzxFrqYpWoOyImuZNPNk2PYjHDeAajmO4er6hRLluXjeMkfqip1
ol57KHzueLlqov1rT3jcNELJAPTYUaE67uj+mhxKyBKkpWyFCGX4/GYI5ixNkgQa
uQpRwnxxFzvZuo7gPQzcWoCds1D1kDIDMk3yoNQ62T6VqGX8fRJBwnQtnfXXBt+S
Nd/oHMk8UY25FrPJbOdsBVjdiEq/vxftfbkISkduINEMsQZsX/TwtzdFfJENdiU5
9dPIXUqlnplSkRihpRQYoCWD2KAcynJXls/MhT5nllHp+wdqyV90qSCeCHlfRie0
c2XRKIzH6VpVGggwFeiZiuw04G5v/d14Za2f3zJ5JxqMAiOv+2LFkjxKb3TBZqPd
wqO+fBr5Ox+zdH/k3qKeMPFuYeoo46l6GzyIZKcefdgjEEId1pVXlaBVt53jlRmT
/Ka5Z6sTwWVft3VhihSiwbYzeThzGf9oPKfbGxAC3EAFS5mSbA1L76NUiLXKA8oW
tAdf79Hy34wrprUjhuh0pTsL9AxUF01Famks1IXBligVL+Ze0MdAHpwcnTjvgLNG
Qt/MFGOQ1otVEPkmjF7WbhkKyCyv0MXd7sq6QJaIQZ30Oz3hzH9KWIeJ8epj7fHR
Uo++27X+skAGchTijpryjnd7uWawkI+dZgxrIoJRiVS/7IRccFQNAPNtku1Nlz2V
dSh7MXZIwZqLqzak+1wwFeKgcME3OyrhGlSJIOhefg48COkWUcrTeNVi88E11pJl
bS3br7e7HonC4+FLFWdYjvotv/78ZKa7pvQxQ2DncmEqaBRWwK/HIB5T6VieX8G2
TrNlLyI0Ul9uiXJ1gj43nhTtjt2u5MdzFaxKpHnS/1Pzqr1f8fJ5W9JIZXbgqm92
1ydFSL34VYLeaqeRpFyAgD+99crd586Ayzj2jRzU0fu52rxh/uh3l9QJMBPy0cNe
eD7EZZXq7ljdQxw8vXLzJmgiFOzy/3hKeIBI5cv+k5eYMdH/UcUm+zx1bgkPFrLF
dfsCoS/+iLRC4N/fOHUdcHaKyWhkkic2W4o3jYZQ8DWPo0yJEYqasJKbaQ0VDIxI
/42G8tLXcac0OmUGJVFdQABdp648x+uqwJayW6KFKRPpztOd2V3j1dSKhfI6rz50
W9gFZKp7+IxBNEo83BZXbF0iZikwTwbr2MWehI89eU23bz72is0/E7jGt7uQSy5p
yBC6HNa4olVOeLnG2mRuF6cUz0axDxG1ooc10kEc9kNMzlcREPa2JPRlUekTzNLN
8XlSUia2LGqN+NYXL8ReOwjKjfmXFc4bGnrH4O1kCiSaZVK7NmIfH5uz6SMsgfbx
yr2vYmL6MvTCLxhIX3l8lEIjWF6G6fsP7JEcxCS05diPl/8+5yQcJez5Ix2b4Qh7
o6BNz9txsgqTTOuBdg/LNDq4NRFih0/I/MErhoeD2cwE2r9mWQSIgcm4nchC3GcS
65k/eEU7lll7Ya3WXVD6eO7RWb9yx7nkbgAzgOjr9hOqc8yXRbbzLUTCwzdjiiWg
TKJlzv9vflFL3cdfgmn/Ed8bxDbMR1FKwofVGkXBW91zD0omfVfCOc6/YveEMAU5
JK9QKBAMJ24UXusi7UT5xjBqFeZ57LIdBi1+LLq86YK1t6U6FMgCzMiKZnW10YYo
+5bSJO0K3zeNRjsUmm4PzhPT+ox5MpH/MBRwpufYQeKZNLafUGuvWA3K5xE53Loe
LxljHlSTp786wOj+i3JmWbjefcU9a8wZBJfdIf8YK5awJ1I0Gq1Im2h2evWSb4L3
VwZNN6KDFcjuEFQ3AsFD2zERU5oM5km2IsqvlNjXOFk/9l3TsuoEMIklY1gB/yuv
7ggnmieh/qJ9FNIiXYFDwREUE9nSN3W2zzidJCMPcusp3IZIBrpIfMjWnJk0SN3P
2mSdyGIzTZzQUKkyzRC6anwkBRMYkVfhU5Do1KILJqnnylb/a425bn9Q4ANw3gvv
brUGc3s/tRyuTKAGo0dyDgXBxOErI6lxG95kM6y2hHeUEgDecWpL1ZX8eKXQZG65
UQ+vuRYMwVW0DkgnsaM7cxizz3Tg1SZorjCH9aU4wtzv6qG4YIjCrjAJ4tu6W5Jx
aAwEdAaJCJHRIVMZZttLGlJOWNxTvCo4Br0OSo0hXc07oOtr3yZAIvzq1LgIrz1g
hwUe1k4HnZqyhPnVoTvNPPi6IZO4TbY9csk9S7fjj16nbyY1iilAZYE9HqBU1zov
YdZLGtS6t/yigWsmoKHDoHfWX0ZIg7O89QUQttLcqoUwmapCAI9iwcHYLec/r3fX
jKIsWMwoAgJuysYiG2zg3e/Mwf+orXu6c8qQPT92btyEfMJJMPcYqnKP7+H2iJAd
JgJ8YHRQVpqe6ZpYTjQYCP3cuxunsdyzhGKLVNUNWe2EwOa7uIgVTOqW+ybGL89A
P5f2ERizghM2iprpd/nj404oful6y01kpxrjdLsUAh+x0l8viBUewTuz2mfIBPxT
ZB7kb2rzw0JK3nkGXRyBt5RIEu3fvoEqMwQZf349Uhq/YNya4rgQEqi7CCgSykyM
/Y0j80xvUaeziecA/k/9/iLozqGWWfje2oMBYhGDo2PlFgzH5Kclr5/U52eaWDBE
SNxmbR5aokPOKHeYDg1J0+c2iJAZuOqwxSAQTc1tVkp6p+hfAUUjAFBBfLCxihSq
PCTj1oOIG98ktijGTTQiKhuL9ko276Lv4c5Sji70LHQynuwKc3serX1H5Y2zNyWq
GpuvOz/b2ajhCyBM3H1GwKjM/ppGtKdWUtbhFAEPjri+RWyUOaWtEBE1Zyj9GkGd
+ME5hW9HLIZt2sxReiGW+Zsj9eT/fWsQ+G0aUa3fgpusTxxdT1357wrTQ44C7rkl
EHv/mUfdkQfpk0BK1tqIfHMi/3aCyvcg1CuFV7o5c0U5EFnbwcvJC/JV/W485k5s
51lTeqt+vc2S1yjSz1UgeoQgoDVjGPINqJDrX3J7e7x+a2T23kJamwA2gBMUGW+Y
LV1i+n67vDn7wyYhaLhLEERr8lvByAcssbWJ9Dz67DuRXi9sehrv2p+1JsH/OmmV
N5nHLdMk/5j8N+3kZR3sVFbBPKo3xMJj9J235IlI05/ls00efrqAyNe8HHvNSmrL
Umcnh9azZMGIkWdSGyz4MCe01vignAJO7y/3L0qYnkSOWyVh6kz9zWNjri0Xod5T
R/V8c3uw4irhj6S7223R1odWHmwTTfVXf/K7lyoPog3wcCj5DSD31Bw1Cs6guNld
jL8IL1d4G4TZwBlKJF7MuLLlLt1gwibfJkg4c+UWoPUq8XR3WjOOJaNq9VXrgNfR
aR+Hbe6AmEpEKu2phgrxbjGPuLzng52MJmUo3yjlZ4Q/tr3y08ePklnhMajAzATn
J82V3ERFU9lWIhvSmZhrltVfTCGfZxAB8tayL7I63m842bpxw0FwLuZuEgcDHoEm
10GZaCV93i8PP32bBaNIx4xA0LIYwC2uTeOQgyEZqPLtzvSioOHB3ImgNu8lx7En
Fhhhnxasyu4J5qRxUMIl1klWsAcJgrdD9ii9YR64YOYgkXFV2hNYCtWfFUao30wn
IuTzhVA9QU6h1Z3bGI/O0KNbrphV0H+F2+EDMIvmzmaTJ0UY6Eww34ZQAwTMRH8H
wwv1oTbRgK+iEulIV/zJGo8XgTtwRMweT1oY/mHtZ3DPiLPlB6NenYEB0svCNBkq
Qc0IrWiSDU2h4daGXjCsprZeNdKaEHEzLnwaT/ggBbPBIaD07ucrWs03Zpp4Q10E
dmI7Pr5+cK19Qr7OYwc6VBXFn1oRU/T3L3jGm1W9E7hEuvvDGiMzSgG3jiDkVdYO
6b+Ywop2OoSBmh1raec/KPnfthnnr3JRp78z6lrvgYdMOmdz+g+Fx8VYL+CM3B7P
k1bu23A2zS1tDXEwxLLd4JcUBosvKrF8QehfQwIayfXnwGc4bleMbbpkGhNcZeks
aV9NND2QWOuZaQjkLDxLSoaG0b9vLDWA0dGbLVGGzXaeosMiQXIVvFgtwkqViRqh
a54V+1nuv2MLdKuzQli6HVeRRSYWhJj2z0vHptchYpBg36LfnoRA7ylVV6S75DFS
kKzTTfIVHVkZ70HrPLqIB94Rh7C5OH3UGPQt2r9ndDEcBqOd8n5s/cE/hAZWPDjF
v9aVv0/YKftUnXPW8XptsPxq4JS7DPTG8Jl4oBuU6/6rMnr+YzwSPzzUrmPg8ISv
MoLWQjx4HADz1GpWGnlluJwoIaoRsz4JXRagoA1JwskCjYA6pAXttDebWSGliPi9
iLLyld0OioJceHJGnrvgNiCsmZZdykpL/IXX/m7L1JohyoSfJJghj69eVCqu8KPv
AZBoMI/M0jpwDOi2yEiHUK7wGbpZ63eCfuPSQ74aHGVJl++KIQGupZlSUFfnsAYU
kG344cxuRzzHTu3m0px3L5+d51d0jVn7v7usH7M4l7nqrTgOqwWfaYQD6BSfEHAN
fQ9hrbO2NLtGSfDBByc2c3MEaMahaiZ0WQ/PDRkyD3d0ILAs5Pb8MePiWWeJj4zu
yKwlHZ7kSr/lbvwZ4idLBpDVNxo5+3Yex/NGp7qz61A4y9LtjrkfhK/SIqUYV2O+
X4qs0T7LA0f29tzNZ9T9SHRyap1DjUb9ZX4CLJkppEd7Zsl9ujeX2uBm2dvZ+Jgp
6/NT7qezM4RArRq9NBGtforHr5JLAEeYQ2PWnORz8+B03Dfs6EYvTcPxsJIwDp/I
7+roOohFAjonI8zLV++RvP9E+wsSohqCu9eHloRFF6oJIt163Tegh8UpfV+Tgx3P
qBwG3pLcDek+dMXmpaRz7WXZ4zqY9gt1LO9ENJZRCn8SZxpX6tA/344OIyHiCVwe
b7gv2dSwcYEfVPKVQwwwvgWcARtxDGsfDZbt/Y8rpm4dC7b4+hwt2KAS//nrMXZ1
hrtPkEvkd/Cy5b9GW/DOpG2HDQzq04UpCM8cb25reaeu9E+RT1M8Jbx6AT2d7RI3
DLcVLJyguEYP9TLGLDPFP10Xp1wReNY1JIm3hNk/BJAUN49PHMmpYsSUFn8DYMNl
iomZtn0jErdE4dZrhbGWoFzplWOToPOirRji4H8Q5b0pcJB69NZ9o9PNJel/7T0J
q6lzKhMC2bfGKfPh06XV5VnAD/Nh4VpE1htQbnv+nd9ZdFdCTwn4jdhTGLtwA7cG
/t42MONcVHa9bNdCdIV77duHWRcZStgdvfBuCEoxh0SUC0BsyRKFtM+Hmjc3In6G
PBRtJ7+aR04bmkU/jsB8QF89JQ8ZQ685vyyaR/nPizn4JK13ErVsikh5rL5aI9CB
mD9UCnRE2n97TSdGyG2+7e0PBoci+IWYc90+S9r+PrGn5CeQKFdYejzxV2IOmait
DD0SZ9jnqSQPeYKaZCrmySRSbD/EQjrxUv+7vDavpQDybLxf2HFxZHNYjDIZrZJf
GAdtSN/eNUjV222z+D8ntv6/YYgyWVys6b+mCRCNFt5xS9x0f47uwyJM2hCEYLie
WKnTbjoKTdizSzwzkSBTOlggfy6Dk8DzObpTO6n+9WjhfB4KX/iKXeKhR7JHHNMQ
C2NfEeKpmneU4I3X6p9gOjxRmQTSOJEt960z3NEC1c8zlJqxDPTE3ieqloO+hLjJ
K4xuJcN0Z4lTEy0SHctKpErHJUPNRIKQqSdF3sC5NsePjhlTBXFS9oyZLaR/eZLf
vkYE8GN3zjnCuqpdAvJ8i4jyPu7BTMf1iHyTElVrqEVGRI0mnXZ/ec+uxjU46sZ4
IuEmehKDyBSOWyasoNuLNj3VTSdoyCJfnx8OJTNaoZlKKII2HezAQSdYIfLHk2dP
g4z4z/s2tesHVroCnsYUNHixiQ9TNePEKUTrsL6DIxxceZTyFYKfq2TU2oroKm43
HbE++ij4qlV5BnbkJ9FN042ugHLOxwW/s4B1xoV1CzIKTO+6k2AYqr2KE4fFpI28
f0fTtlVX1YHsG43JGkAwQ8jmUoCT/qgS0aMgx1OzKjDgY/6/AG7q8lPjHiA8SdDI
y3fFOs9BMAzEigZ5ocMmTl7hVhmGAptRGqadcImh4gKrPtnic1UWHx7SFjdasxqA
02Ef8PAY9ogNjX5zK2diu9BKjtWyF69XBkgxsA56PfVhQu6mTViPO/OK5iGbNT0o
r1Dwx3mStUk6W9wio1M7V737yoCg1o1eQOKg1diBRm2WMa2Lbgfnd139WGDveM5h
cfYu2LE/VBu7RDQCRRwdyooHGT/WlH9hujFegSne/pvBRQ8L+pBptwzyniuT7Vay
AeU+4mKJ8a0Ejydz9u1iixp5ZslmEdz3N8YSzpNQRUhEKaOnHZA0jMiJoFt0ipaR
wSRShbIhcn/3XeeaYq2youKag/9PZvIw2FcW3R+bxaEsyol/u8CshsKjiyjQBldN
s7guTdiwU3+Y8+ZgZ98G7m62yLZYEH/Bf73UgB2Mne/0P7eYJcuFnhfnJrqQREbv
HGqID61VLaaigHCx8l/tAcykJaaH5PKDqUJF4o0Oupepdn3ZmMu3TXsEAPgm0hjD
IyNQvkcYJGbabDzEKnb7zaG7XkjlA5bwd00KBRKQ8/id+wAiKdtkiPsphK1btDMm
rbTbSJe65voabnQ5ZBMxEoLaciiTN3Ot5oI8+kONmEHG1DRe8IF/gmaWQq+eFJbY
N+RU1KpSlOeXaLfqXKc9/jZoBdoEZMnHU+5cddC3LWuHsR2FIWBSV6qmXKkHsEr5
2ZJ+z/zgowjC+wF507W8dFeA9uswzpOP4GsxMpdx8dBAv37BgderFbjh4a6ryfy1
Onhp9Edg1aMND6+K3iGf85AfcBybnzwS9KNLAA9lGfdFqa4WZQpNUvIBY2/BFFqx
xjJKWk7tGaK81vu1MefGme9tP/oFlTTWi01LLbJ8ififFDLRwfl1CEw7L2g5l9Yi
73GC3UMPJUl1f/aWk/30q+wLNZumx2zuPaBVudy1xCM+askmK1W6lcF5kTrELzre
HtYDtD2oifeI2McNshtCsKLtE0cPxn1AqkPZw+aMznydZqzRHcSPnURAL/RZNMdo
hOfcTzEybRj/gOz20YWvDPqovwuro2HlGuq+6EEHgiZ4stqUue0CxiKZxNL8gZcC
Fne08OfyXrS7h2wf0FPFzy7sANx/Lp1e3OGUQ8RpNXjvmTCyNf9mwHwQILIfu/Ax
SAArFlQrgCqh2/s10fIXqS+lRQiXjHsweusDQF2MfT8TvZw5BIi+3M8Tj4+FoW0Y
DMm8/PqAB9o53gwiIJ6qIjev7mJpJwXJh8QIbfGXS9+eFq9AVbFd44u9DNIs14Ty
58yAvzcXPjvoTvlaV5ti171bxE+y7Lolly10kPNJbyHrVGLRXx8uh9aILvE8yz7Y
haVW/ITFOkVunds+M7BFzbMEE4B9Vj1fVUy3SjcEww7VUyHcbFc0ZPBdT4WpBWUl
Ljlz/gcJRYbOpa4Ojgatktsz3aCPuLQLg12ivGyPrFPcD4XWGf/POqDCZ3Uy5oXn
rgmEAyYsibVHv5LtQVWg4vdG4oRrp/F8P/OABkboOjC5X5UkbnujWjjisGyzyhzj
9VJSMn68h9xjxDnEr7mpOSuNei+do/GZfinzhyqIayOhqeEzwpaAiLqsv4os5iys
dIF+N7hIcAi+oyEw4PGyHydC4QSuVf9cfXX+geNMOM/FoMAu1gGDda3aEi8dNVOm
Gv850eAvFUz84H68nkhc2A6a6Fd2PCcJjqewgTbwAMTT/yrtHUqFXhrqp0yX5vcw
73P+I9t9iBlP++Qi51chhqJZN0wYWU1/Fu0SPmgglMYYX2rEUA8IrUkPwsHPDIcR
WbStfcfxABMEr6WkNL6X4yvWaUpQFVlQxXLN9OdhojZ7u5I7osIvliyqXXTH7aFh
4RxuG6/zk/DndyZ6GeCHkgpn8I6wOKKVzJx/dlcL1l1lNonb00YUNR1J8nTdMCN0
wqIXTAOyRRmRoTBzmp0K6PDZOSHupMi63hUTyymlR1TL5gKQ0wTyOnfJKV/A8pRH
cWaFaD0QIJv79tRhPbJFZqlC9Q1y/WhvMCwxZZ2Ma3rXx7FQTjOGh6ReQMLLRYpR
Iy4tvq2FwTgdzFZsDPHnyhZSnkyJqeL/D7CeGR6IGOs8WDlQx5hTz35xzju9Yfdy
FvFQpA3s2yeC0RkLpE+v4BOcfSHSJ4HMYbITac2XqMdXn6ZLqVCXPqtJ5FTiyH8v
8uYdF3dzW5k5jXMPaUfQvVhvTeceq5dLQRFoo10gLEFWfVaoixAqFuQLf7wRhaoO
KLL30ka/inO9uX8sLyehXoV33+yfsSBLysZtmMZ/5BOuGZUmYUhD2dbiJqMlp/8o
bUJ9XR6h3eaM2PIfDy2NFBUXcl4dfgFRKyXSiWiX48J3nCdshBp0JL73UugtSwkv
iXku9x/y7LB5YBHUVzqDmCr8XmcEhNb/0Vqr9PGoIf8lI2m/9yVFXPjXlxjQHhKp
UF+C4cXeJINNo3Zel0rCHjdifH+242lOJSHfBsZyedUr6zHV5fj32l0mhzwpFfgX
m5HR2lJ8Yu8inpa61Yti7lHk1uu5nQSFQNL0F07dsYQMnkNceGu6L3mWsOGlSk0/
o2ABJ+ErfhL6M6uH1Vbc0Hd7fi++E92O/uSiOViMp8uFUrkSKb7B88FlZgJ/s1KA
AXbgFXfFYChZO/5gy5+kUPvCO0wD1+8l2atXI/c2g/Of6agj79AOF5wC2xx8yiz5
4iM968blVd14gtTxJhpCa6gLNJQcecDlar1grPC+bYnqHfKQVTgNlq/tPKh2WP2t
NtzUq3ux1EZYCRVKf7MC4G+DJk3HomFSUXCNqn3laYuS4aNt2WCBeUv4HaXEKevQ
5np16+dmFCWdugw3Mpa2/7DSX5qO+0Mimj53YqYty1b/MRywJXpRhqJZI//lnj7W
smLV7qDWGq37+fKTEK42ynSLOlmLNLMbX0MB4XV1BM47FPDmFfhPLPWg0IzmLgAf
HJBGTxMqGuowLOERUq7I3Ua6meT1zZGcqHjBbbE34P7Exby4Q4Zn6RKQP4idaERQ
rTvozuQfCeWbHRdAxnZfRTsjt374zYLhI52PX8kbEnAl0SKTrvtI8Ah2QgkCH8Vq
I3amJ0IAzDMDjRJgMJA4nIftMpAFzb/Go0NPEH5Pon9iwkhUvSE6ZUeU+L7961xA
iQz2rOrp6oiKxgq8qFdL/iqoRi3+MnWGmiggNBc9pZeoXdvtHjxmjbGvtocdLas2
L5JzzfPPjqTBJSVBt0jTnBB8TkP+gnHZNcMlou2H/SYR5OdiJyVG4iRbQGe9DhgI
Nnd6KEm2RpYzRGgTYQtQITHXK9MHXFam7l9rlYc6kwTkIkZ/myzHS/wg70EmE34v
yXGgISg/WKxdXv5N0vXcpr0ddGjS//yguFWCv0hGPLbxElvHsYCZdmdSwzx002wH
gEXlUb3U3XhG/nCkz8sunrKerZlQ5DTb9tLdaiTlQbEHqhhs9jaFutTENHwGrpA8
kEwZ2g3rPcZjt0V5INadsrrMFeAM87BeSeAeRZiAPxwyGVBdFPYkhR1j3APpvQq8
G9qeIXO0Wy3eMrT+jB+33Q/u4U8KjFKuHt/zNZfmy+K0c53XzwBq6CScX9lgugAr
Dwu3CJ8TK4taAtSbCFdCFysZAbvskph/VlviKYuVq4GQ5W4GlnY4vOHtv3wXzrvc
U47+sWgPCzzdKhMpj5IyKSljWYNUqme4/PGgrKgCV8w9zmgnchXLeb6l76HwIg1X
I1LK2C9J2ZtZwY8moRx9K/DlpoGU6Od/SRF77xVw2ocH5adhO52F0ODnuABfqBaX
g3W5aSt5uYrpclGysY7R3+k8L77XTmvpVTW8Dq+hwSb7ef3lY2HZ0exygfPqybBq
zlxprOfjrocj2mCAB3pIZWyWUakpZZN+u4dFuLfDISZSY10gcLh/U3RlhEjMVUbz
JIJxKaO4eM+Xy1paMshxdOI8d8pxywpJ7x1e1xwASD/BVuuADB91h/mG4/2hyyKa
l6QXQUxayghgobeAUKMva2frxTtGMgys5ASwjIHglyUjmAWoXUFxlfSuQP8FceYa
F8jtbju/I/mtna6kCnfs2cCwPVmNGRSf4T3mcgFRRRLegbbogDTLZu7XnFFBrxiG
YK0+ro/diJZL/tGIsqH4B6XYIP+Y1J0oS8lUCXOyk74sqpUTvRSaWmAcBCbM8j3Y
/Zw+5tuqCn0/XHHjVdR73R4gvNqTW2gfRpMKPYJNAZdco6QtENeBJuU67tua56K4
l+yvgTjlY7GbsrnxtyVasDesk7cn53cKz6F63plXQz6XZbBMb57YrS0Z+d4vuadi
R3jEa2kLRKsyL6lfApQdAMzaSlcOc9m/MATqiRimgC9HuxyvG7M2p5TLozKGGLZj
sl44+qRSUwF7lMgi51kEMPPDR9nXa71EofbIDazm7MqC5gwClOQPibtCZ+lZUsQ7
M3UTWUGiYQl00eTDqQ2vsNdds/jhf1LO86OuvJ7hfWHR/EgPD8OKV1JL7GA2BdEP
hPZ0dkkiDyHQkRgoB4XB5HxCjScYiS9dxT3TY9EfyZ44JCsDQF2D9Uc9zJyA2dk5
VZ1zIp0MYZ2gVgiGnkJVJsiYy22baVl11uC1P8f+n0zsrPx+ODyO40NthsYNcdEp
Xfgk6UevmEAtQa8ePfWLmmJgRvJbwj43MJAqyMBVZIARY7kMobsbrbSdtQP9Ueof
fPquWzP4MY2RIAO8uXWohNdCL94PQ00Yv4h2cpN6miwCmTWwc/BLMrI9zPg7Ni7B
iTLWByUeT6wPFZbIi+FdjCwuKqYbMDt2uT2HDiGhNO2BSDj06n8kgTWuQahihy++
2JwcMSPYUpOl9my6BJg6zM1kXljDgGYqMWIU8TMfZXOOaRiQ6kLLlK7NQVvv0s1p
fgWWov8ytlZb52mOlLhX3yR2ZeA4M9QsHG8urms9lYq7Aje0HbpCUOwa1o/rmYbG
I5FA1VER9QSoSpgr9Qe/GR129S4AHzbcEDvW3A8g/Rm+6QMnwUalblDPFAkdlrs7
SZzcdCLLvAt6FkLEia57y5XyoUznkgCEm3hZtLbviU7OjIr1hZzaQ2GSijat8u7c
m2OTw7iJwXfjuGv+aavcghmq3g8ALHQlRXlprVeiuv1+lgUn8QuTCb9E3BYWi7S/
g1KHan0ib2ewp1FBPU7wiMPE0ySzzKUSns92ZziIUHh+tI90Pc6AEng3vdL/B2A8
WjhONn9c9BoV0VoYEOVztV1Z+kXX+cYCZ7ac/CMMOxoSfISs0LRuJWGVQVbO6C82
jgwFj6ocNYRC6ZmrhfRTheliGsCS38ggOwgAu+/sL+0L0UQtXsTwbMRL54K7hOrn
uAn0u4dCjkUmdIHvKkyGgfVxVP4wTLVCT0FcY0O+9lJayNE25hoOnS709ubPGILc
bykPUDNE2fS3MkGw1NoRRA1/tXUF+WkXKSQHKqg11vxwC+uzGE8QgEF7tcTNJ/6C
uu06KCp5lL5wL9qk00YgSSwnQs0zN3GjLHU+e0CWgxW/6ssu84LJbTvHZW8rpnPQ
3x0hTj7WoqAOwvHlcqFZBrYXw8P47ORBcWjYXErJDqEfoxVMVl/TkECeITCpK93L
aN3DOUXikPDtw3rJFoMtd6CydUCGSNQA5Fmg3+bLtyZouGxI3H7gTVlUyjv3mIJI
sCzDg7Rc6ZJIIBug/+bbHpJaCAwM5Z+KAZp+QHQJdWjgksiwHJG8Vste4Wz+sBII
i0APyzqeTYwjyc2uEQr1whRh19AiVkKhN96G//CYCxAMoNGg6Imt5N/CVYsoiK/+
xL+SoXWY6KZcxz9xU4K/NlCTvSAurK27ixKDI8MKR9kKauPZ/Pne/Mz3qqyGP3YQ
4T9vR3G/4341Z4tCmE0trYu8VxsZjKEX/7rELgSS90H3QZx0l4tnTe3J7TfSn0dC
w0TVHqoy1LDhIzpPoCWf3HkqXP9OUJg0j4OygkZqXgTXV3Q94UZK1mv8ptcdGWmA
PgBvIgFeWudkzcRfte8AXzzihXzQiqC6baKGbQlXTr+d22kEH7OhjgJNKolwjZdN
vBMRQviCklWqpwmf9NeAj9IUziyPBBkyIHCWOOUtqd9vooYCAu2eYad3+YM+OyU7
cXr5O76ZZO5T46lvYzvBHYm9xSJSiNNbDNppOONYOyda7JHJQFNRMXpIyJyH9fXV
pGcAcDEGxHViuR2Y5pQA4o4jh1zabhhl3tcJogIdfDPMvW16jkDyFalj9yWltYvD
jGCBtGpldmO5y9kUDh/oyTrksk9a5cxB+ggp8kJELpCfyGAjDJenkuW9BOBlm2Uj
0J//VjTQISKNcUeLI5LwurXSMbZe4Oe4QFj4RFMrXViSIRprgnT7BUNPVSu99kWE
Vu/FelpAD1Z+L7nrgQf+8fz7nsICXERapERhsaEhfij9chq+wNDcRkiIFOrcjgN/
cOH1gmSxxi8ksRXhN4PcpiPOht4wszTDXUa4LBCA1SYjRA1cGdaDGxHIQH4ncqmM
ayt/txdoFF7CPOo/4y61miQAbHpDuQ+gGjtfZcqOEBeXrKJ5CoAydF+LUu29Qqkk
ElTUxkhed49RaUgoX3RVG0P1tn4ep0T80ohhZqJl5i9jygwGbo4h8Ug6IXkrnKRH
1k8e8VT+/ByWu/IuwaFWxvBSvDrhV9RAJQG/CrBmvIH1jRwd3edXNNf18Z08K7bf
aMOkdAyOVEQmCRzADG27DH0fx06Phg++olAQyJ4ICtrK0oLhegLaisWZ6v0FN7YY
mj5aJQlaEQ54gsodMcW+EwEpHK/mI9JLapWqeaWdVy2S949vSFS6O87iEtNZ+mTs
/jWy2ST3rJTcaTRz7BO07CeVIsS9O4Gdktaz0OkyUdqoEnVois2scLY7kSNVF6Un
GTaDEXug+zqh/cLArtyBV2lJThZQaMtmAzjKUYOMO+8Hey5zeUsy4LiijAycmsl4
8GZbXCokFKYDWMQvGRCqfI3t3PFWBe8m2JMim6w9+M3lniZPVsGBSVzF0/6/ra6D
FhbQVM3DUi93vca9P6lV09WyhEErCg5cSNXRg3wGrQKP/PuZMwtEOqxB6i7hZ5Ew
dM5bEY+4CEHJPjCLNu0FV1E+Ub+xwZAh0MdX5Vew/ICX7WU6LdC4kQWFvKGmVIzs
Ff0ZYklj1Aphaxhkw5BHRDDtq7IHvV1cAf3l6DZYliSHGPBpgaVK13RnEHX8QTjf
Z+zQZek4lm20pEkHXBko0HroZPF/4oRTD/HgvLbm5TxOCUQKvHVxboUNSijCkVUt
bsuc1W2c1TBtSNjH8+zXTqZOmaAIMP8vn8xbLiOCjpfWqhTctQ6y9/6OQvfYLdSE
VNCyv3sybVVAo+MflHcW8WgBBb5m4Xu+USSqxD0PowjgJMWFNlj/D1/jAPYtTvaH
bqfRKySHtPMh5tmQz6AkWbQp+FUNMWgeRPX8uEW3kJaKN1ZsgruDySQ0S7+dgkTM
lfJEubdrtU1Jvx9AnAdvKD5rqTddXmqWN7ysh5aHuSgaAKj70mFkJ1dM3ZijDOnI
TEjRI12cC6Z8oUOUvEpT/xHTIez5s4nxndfsDMyXAFoEmb8IAXqDbSJU2dFwebYy
H+/3bMG0ESLgVmCraOe2NCQ+ALyKJcMusFJJ4cOKJ8sDZ0zyyaCf26FM6t173iRD
cq7miGSEw2x5zm1sH6icPFHznGYXQrzHkRCwAPgRoZVo6VUWvCkit3k55M2bUqon
yCMU5PO03wsxPiF5eQiqjIobfeppL+JUgqPDRP2v5S2pb4px8cXuItfY9uLKq1kE
Cy1LelnSKPidmT87e/6eeTyVrbG7nnQ5hvrlOwVRe+ZHxQrhbl//wuvYtlmJEgNA
+7bajb3FEi4pavGRodRV8OxaEIui9I30Uj9RjkHr0wxbm0JwvpmB8BKW9Q2yMMqT
aTD0VgocvWgTf7a4JQikaiUmQoRPWIHMRnrRJ5CbZPShJAWxU1tx7R2wglvxmLKj
9fZNjt7seKv2T+/GP+FyQKRi3PjIf1KsSo+GKhHwBXTin6/hI0UmkSHKvrwbgRjk
hTtNSwJ+aMF0RrrMV3KmFM30HxC5bxJ8ErEYYSASOmXbKjVU6E9IJK3gygs6igy2
vU0oOjqxxJm40rv0n8PYHct/dQpvwOFHPqUwKPt8sN7mzKPreT2aMlX5eWciz3nd
u7c38H6uu8xQB+7cTAl6YGe/H5N4LdlIV/M5fsb5obiJbD9NVZShApZ14qb0odru
5gMj8TNmgHyug0AtVsnAxV733uhXN1yc1I/lk6tWv1+SSjlOUJljgJc6CQhhOaHq
vr3X1ckqqP/sNd4lqWRlKA906/aY3J8ITBsRcLsE5HsCHyzo9QTTzaZz1YENyjDV
`pragma protect end_protected
