// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
DSgsJ4ZdrGY/yR+bZmUfCLH0rmxLa/Qx1pSvYbu86WY3jlI3hgiCbaMuhTA1LaVd1a+6HWfQIl07
bbPM31N4N5Q9aIgVBCEV4HVDmK/vIp2CeZmk/1IR24whRXqXp5FjqhkBbYGZ8uIJOb1oP9detv5W
c5XOt6tjP9g9sjUd8DfFCybsRMYcXm1zFtaf0o3v4B33aNPcPv6JKtdu0NchQquEPP1wa68993NS
GmuVnN7Bwj5wUGWnpG1peIpYy3+NCLqmnddIB0zrNtegr+vm838yt/y7Q6xjMmnLqiD6gCSkNCQv
y8Uyo9gBxyxuWqulXKq4ld7xoYWYKEt/XePDSQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
rij6LH+gA16MFCpt7jCg1/Oz4s28Oyn4iBGv1I1HfEP7eh6WL9oPPGIFqMkl1xGlRKwx65XDIYL5
V11LwD1sQysezo+03PxurF5xObCpiXW9kJrLXG5wWY5JH+JWx4wwPGl+NRyJDBSZ6EJ+JEjiDUiQ
e4tXxVYaBgz1ft3ToDRWVXlMGWzHkEGO6Cvp2k4z8Y+MKpWTdvDnGEDIq0hpxBaDRASV5WYuEqlO
tm70P8NWoYHRSWlxRewkCokEkwfr/ygExW+1NdLdv0ZNySAIRM/wBoOeHzOVQ8JwnOTsI8puAbN3
AZrwgjsUDlOVsSVBk5JVkZr6JIirWaqF+4E8/FVWtE/ocBkfyry7UP6zsdyyySRCOaNR6ic6pxrl
JQP57WgavR+xdUhq1VUXJqiq0hqKDwkhyQ2cBolX8lcw2PmicpM2TnHrvQPbirLyAUKoEpZE4zT4
gBstMu3W9m22vWsHlFxPofTCBhKQwPV8vUkKvJ2VNgN9vAUxTOtVt5HYYQPpzQPJfKNLtD8DBlfA
avEFBdHXSAJ8MpOYN+Gp4qz+JATjwjn3mp5iaTgZIOjNyMxLgc86dKUC+sVPQoaKY7V11tFVFO0f
nnknL2phFXea4C8WRiWtRz2ymIi5iuHV5Ox6r30iqyRTregHuPKr7irm1zOWaObOaHBqZmSX9SJZ
Fq0acmd/nX20mZVsJWr8RydWoufAGQyeCnsQ1+n/d7mVEEvhFzVGrx9DI/iQ1OR3lPSUIkApAQUt
ko3gc9nlpCXCQuOMkeDroN4SIP97ENJrBoLUXVl0ic4ONfVfpSzOv3OOpBkyaqJt08avlfj1o3/f
ACyA6v5pLEBUr1PDdxirBiVj022xxlAG+8DTwfmuI5aC3roMKMvDYiD/ZQejnmB2mkLC3LKP5eGk
ArIix9l1gfUh+quFu1Gy04Gp8FeoY/B9N6pbq6z38oTQUKicnqm62gZUHrBjsLo5ge3Bl06J2ugj
Ouu4bR6gLW0z4b0CNcKkrNB99X2VPrct/pagxlpKSjn4x89QI9fa50y0bTzRN+U4N8W88bfwfSik
uqAIdnp7zVij/5fplMX9GoDcYA/kiMJ9f9/+SzbDH1rOJZaoptCckBpGccEahOMknWsPDXxgjfmD
H2/S9kxEwrcuZ3Eo+XM9qbLCru6SapHMdJcFYDsGRX1UTjsMcrEDv1s+PAmb0sYprjgK2Uin9ffW
o/Dd8MSBnR/cziCO1VQ/tNV4UiY3fdnYpPXcpz1RRVAOzLxss6BlJRglxHpJ6SZJV8EuE3etgVk/
eWHrCc7wm5wxNRj4Mn+sFK4Mqk0wdXOmebo+cVGckpytYFMcOmRnF0PzAuXek76qt7BX+z6vO645
g4AfwjzfkUJTl6dlI0vSVnCmZn1vHFzzxR7nYEO2GCpr8TJwh2hYzjvGFXdgvI1Kqt3VrjqFhz0l
XNE6AAxcvFjzZM8Zx73TnxRP4veFGoR1u+AsJ0OHZALKvz/BFNqFFvLjBhTGogFbMA4jB5VHS0QZ
HotoKncmqCgKk908+UCw4xz9rhEoWH87qP4DdVZrgUuTEvi6GxEMa/FkFKHlZPsRIOE6OM8IGgDn
MYG4X8vhyPZI21dNmq/t2xoUPrcwWsgLWjnv49M2gR7kVToXO1GEEdUzt+rqZnisKqtxvyd7VLrv
/NR3SjoD0HO8LGU4dHdJ40jK4I4Cov5TR9uLDlbRppCRlxuPoLeYZvD1lbWTR7ugcEU9LckUr+x4
yXORahUlvoqBH9WNSUUH2rpKVvdTFZmTUOBTRrtR+5Jzfo6KLmmbdMIXJKYm/tAro63d1RsSqaC9
e74frYMkVfnpzEHl1ZcQOybncfNlSW8Vc7XEmW/488h6BmgR3wQXELywFdVYiWvcx46wfYS2s+4f
FVFO3LlJEmB2tChBAHfC75N2vAXCBjUj1iFweUd4CdeF1rD/8BWcpnMkCBWJSbR7k0qCyzldTH9v
Qp1KUrqIcwlMzysDFKF9JQo9kKgybmgEPB0l8F//gK7YH0AkDFpMj9TiCu32BIZ0kGHcVpL9ulaX
6Hn3Gc51MJMkCSTAmgh56e+PBJmZKBd1/z0SsmmZ4OOK9vHwzpoeshapLLT6PvZjh0wuEjGVUPQx
3TJPMxakuoSsnd/Voc1CiRbdfLZk0dotOFPxUyOEl+eO8aPzhbXekMEVGSiS6kgulKAiCA0sW5tR
GBwo4KXZzNtgG0dZn9Lqd9BhddCku3KO3HFijoJGnOwMMdmSc8Pnz2Gt/zzsKY2YmvjZpB6mYn3J
WmvGixSA8fVBKnGiJ6/B6Ho66cwD5xZF0rMugYT3cpnyoT8qUIFPTMLkOmnpgFbUyVmK9IYuYB24
3EGvwFeLWLahPsKM0tCQy5oFF/msoBZjnL8lfq+r7zgzsMjLKA4Oxk9xVPAmCAjddoHbDBHvoK/C
6YI2AdrZuFHTF0zUJ+pa6L26dCvPntgR/G++oe5R1ueXT+QjQ7tsTQXetT83D4HKJuxSlvbPGPDw
lXh81d5HLueY8lwjeBDAbsRSAMuGDX8dhtinYTnxWwM1Tg21kHYv4zmob+Ld3hxOuVy6FDKKzXII
Tkg+gzq6/87wVV/bEv1WUUWsoVY7W7SFkUJRfQs8uly9Jwgw28S6BD14F1yYaxFizcbtbgXxsyNu
E1Un/IOhz/Az2pCcrDSW6iBLnGd/wg5OeP4VeEtza7DJoypZJfntKFmxJQEDoS3LglDgWjB9CXbJ
xn1zSnbzWQ7HsJk4L1dgfZbrcrRr8YaUapgaOYYwL15bFEbeHmeeB2Wd2EzmbmYc62Rah+JvVUrh
Uizj35UWs+b7uv1kX1S59hkYof5hZy6CB+oxScizAOnxEq2OHBNJsffHecx3EhqGq0jiWaNmAe7Q
bvb7XqEANm+aS7sBM7VnuUmZ7RwMKjyYz1q8JHPiavlAMg2dvH94KdIoNlh05oJZM76Lt4WT35CY
+zErI2Uulf4tjhTOGpAVPLwHy4GcD7vOGIMkfXlDLB4R99IMnEk8FbGwrZ79N1h3cxmfPRyDgvHL
bcaqnzqWY+nW4i1lm524jOYNOn5vkELGAAYZ3VYh1RKk8Yc/OWXgAkUMrCs+kQ5dGDlrQbQGfA5u
rla9syud4MILIjiTnTQnqzF7DM7ObYXCAxmQNlZaCduGnMy4hjV5R0zpOHlenathHeOoM3/2/1j6
gu+AXRzyFJMH5tDdNTMoWThkYy2EfGM9b+fZ/tdUxxkvEhNejeqJS8Am6UpnNeWe9+OIvi7BA1T2
iA4zZr29q8BEQCbdNf9S3QiymDErThGqX5+egWCmaX7mnfWBSKwC05ar0ywpP1bCIwtl1VD+q1gA
ozib4d3OfXxKeLB4dynTlQb+ozYqBYbL08EzhA7kVWbBIHKdIWrEoCbHb9nj52MKFHW6mTd5CBk+
IAk8+9KApeqIBuPfs6fM4uncvtSakJRksqD8gMRSqXHW8u4Qc9CVIGRJGIJGTs8Bg4oIMIFyHilg
o5DHhfbSsqn3/ttoDLpHI5QSCUxT2gRM5z1yOfA80RUkOky7BH9cqS3kwlcckijbhbdZ43yKOHWk
aUG+9cXU3ZuZyqGe0QRaTNRGUu8isxlSuMwlTKuzTKA9T4sYRWfWLJ3qf0ixVSlYJCHoNdd6Db5d
2yVNriocjvt29f79RHCkagiCsbsp9tVSjWGWtbWADocyiWPYZpfJyHGeKCSaeuLnh3Tz6wHcvTX8
GTZRlRsuCJ6dRNqtpgAwiXJqhf+bsY32tR60eZ39E5LrJViXpOtDymb0iIx2pmzZ/I6IgNMpcdhq
YedBVrZo9MBosDC169+FT2PrtVKP0bHVhhAvzmpBREi5lXDgnW59Ymtd6i3nTKerUwV9SjOZOoCJ
EC4GoKMgPjcZEyb6whR+2WGwyr6BJm1IizBHjgJCcGcXqIhdYSx4vl3D3cLOGrNo4M+G21gyuTl2
2gBn1BEkxNIFhmM/ElNY+01jnRK1zUtnOKTLDdJ2apLKlnvLGJvntyKgPpd5baYYQvT5jyDO7m8K
bOw7Fnilof3GOJF40jduc78Q+lfqgzqp27QE14BfIXKdOM8O98/hlxLTtIk+TaUAQ2x090k4Fse+
7oAI6QaRKt4OBDiHLBhKwD5aaJK2rB/a4piSfNfEKfmyd3tnLY4BvA4PDKqbh5H0DKL3R5OEUX2o
DHLeRajyJUK2yNma80hRoOnZCoP/plop1INVhDaW1Y85uMM2jjTMH2BHNN3X0K/IK6/6JM1Xhwh9
jIaaQ+yMW6xAgezCAL7BhVA5b+PPyqWcIoZuzZVM0nrYJquOc8Jr1HS4r/bf1tTvk7/u6Ij3jeEA
oQ5YpSnYs8oZ+UK1szf4hiNzbxtHSZJ9h6cGLpJYsP167a2qoIPpKwaKSXYTYxLfkL7CCyjK05Zv
hpzC3xk6qhe0hqJxHRM9mHkGbern77ExvJOyfXGix8rjBJBx1H4lzSMLfTSZjI2n0elpVlykoeab
J+jPaSO3XpAbuuRl1Ucdtv8vbcQ0HkMxKPf9h7uMMVW9r05Ixok1hHth7KAhgG7+oBwhwtcs3XnV
xXZoJcpJeEP70kt+fX5O68xMVnlBuD0n2mzi7Ko3+nvoQdgwuq77fhvdCEcFYwl2BxcGMS1yKOF5
lfLy9hBY6b5D/EMLy0D1bya03VDofPXPgFnO9fOEnRI/x7RSAv2Z/+ZWtZNzN8axRoSHpquCqXbM
znfiEee0o6XWnO+wcHHfqyY5fV5rTIt2/r9T6Yy59BME6qeuKsS2hxjkm9QvpFJ2S6eQIT3Za3sZ
5C7QruRcduQgF85imuI0Wa9t+dRcuYj+1Kwspun2ogsDDzO5agElMPuev+OeR18WBGDNdvddtiZV
1LiaMt5j4GPMnVYY7Sw2XP/TQOxenVU1JT+O4fEtg/EcSxmsbHbYkTjLFdC+RQNtPYWaZpREMEyU
B5EcORLCdcuCxl54z80qxjBmVp9clseCPIUoRX+MIIFZQ4lgCmVaxODIKkTyMhrA7vkdp3LMzy/M
1rXJ/j34y8L6CFg55ddnYxlI15TciI8Xu5xhMd3CxvJ3Cfzge5eeTy6adp+aKvVAfhUJuYIMnJ2g
/STq6zC1/rFtu/bUTznsMGxp2Wkg/MZH5a1awsG0Nn0W0vEv5g004gQAQJqnoXTBV7w5G46dd84f
S2stxPuEUgHZ9Z8TPjzXs/t1QnxHt/egSj7BNehLQ+gZ1wW3mrHf5JaHoJboiAi1eZT12j3tg5kq
fUdyxwJyr3Gz7HWBCMf6FTEBSGXEfwbThtA8YxDgDyVBjvWw8cWxcqwRcSdwNlvCDZnhzuu9MDVP
aVNN7ivzI7LjM4Q2fUPPMiQS90Gitl10fPVM9rRuHQZF0q6a2FvCbiVi7aOrxIzqKL3B3fsk1tYe
f3R4O91kbO8hEk0u3OU/AM2F52CgrNT+LW3rs5yRiFsS40alcVY/Uo22yvfOg2EGN2Z7imQiz0SC
3U+t2tI3YlHbl47uoWaVME8a1zYJjnJfTBeFiyqM/zP7jClCrRG+j/P5Up/BSsyR6TAmyjI1fXkA
DFeRh6CLVW+LoTC7KrYeWw5HTUptWZuBsN/q6liK1SwCvbIfl1XWEVnVbhWoIB6N+U+DRO5RoYUR
jAG6iuy3sK6Dim5Cjhh77EruzqO76p5dUc1DJuKNRi5CPjLmUwp3aRQHxLiddjwE3BSeV/jnRXha
LXKYsG4nSjXjPM3FA9xuviJYKSS76aIeDPhPRZYESX00XFmwDBB4p70BFvZVZ+a27OsRvn7EjooT
2UWBdvIky2rMqkaRFCKKbf/TEKMSgt8K+DGI5zki6t3PprChDNF4CAFbpzSCDDB7n5pE+ETw0acD
PGgCTTBJPxBG53WqjRHnEx5f2n7bo6a8IXjxoKBx1pJ7CQ1PPDLZQc6jdgjwJxFpLkdJq2WDh0DO
6F6Iv5az6Gmrbhdx92qGqyTUt53aOxPbVFkjMn3/o5Zw1lcSzcYTFVttN+H4ILXb4DCBsSc9G/AH
ba0ORwQkhUwGSSKMMcZIRJC/ov4YvAtze7bjB/p0fPZDyglTINtMJcl/WVIyvFB7cC4otw3Damq5
AqajMmX3wFqLZg8qyF7rInUp5qcMb4RAnmi110R70L1hv15kMn98f/euXnvP3+Td0fexK3sZweKW
1OWNo5PHjOtKE1bVJEYeVHjQgrqEm2RVvmpFP2WWBUIotMMnHm3FGTjkZZpIoyPRS7EFTjpyjO5m
uTfMiHhbIM3y4c1bmMyVsDNwgTarKO/52PgMpajX2IBSPfZAyYHcAYx7Zf+1vSmUKC++9jNkFOFr
8MYGvipAvrp5KpWR8nkFkREtg3T5ewoEGydd/eLV+Lxu99X6KxvNrpQ/QlJd7Bcu6uDYnVWfh4L0
zut1eH6mXkn/9iil3QodV9yGc7a1f00jcyygC7TaDrQRzJCs07J3+4IGPkM/vAnufgTpKSDcZHMP
iW+8A8g2r3FPJC5Uc43Svg4mJX7QaZh0C5v3sNLwbisdf192utDFYZ5IrnC0UAu5mTrIzvxgkzO5
XbcXAEC856AUfIxbOlfO4p5JC80PT1Yv1LfgTESDZ5cslEnzS6nOLkBZ35VkZGhxnxPZ1b5yvS34
sxBJiXgUD/+jM5aRD2nL4HBor9A1UmDlP9OqON8PbQKRUD36kLJ1LVs2XVMqF1Jz9+emebbhq5Tm
ZvWpbo2aHSfYUFDemT5IyULA9FUAEPyJmfFIgI324UyXRPMas1pbWFUueRqx29Dh4NFeNSQrhBc0
hFy/GFoRK9r8ju6OP/a3Nu06dkoYiZwbViyJi7duRkl9Wrora0jUL3mXzguYbQ3LK9+PDengvgKi
mg7WcCnBkgTC/pqCUKXl91hINtlVohhj+SbfhOv37gUOO70bh1VcLyCjyElRi+BDaPHyl8dvKCx4
uXaA+g3H/yt1rpmS9TE8rb9SNWZIbJzYZDP1MO2tOBhuQF4TUISJXIxyJJLTL60r6WpqtNr4d2z2
+VtgU2BB+qfzzuuRLNBMcJZpFtczXIpsJD+mXBhVPwIhuFv704RU4lxEiW7MJ4SoaeyqHKcSeF5e
jXmwjw6fGtRswzldcJQ8y2/o6iCSQogc54hE35enNgCzPVBX84c+HFR2Nq1zFF1YPbdO6ytXcey8
Bw27DPx9pobx5vVdNg6sb+FyWHUYGAUyJugu2AqWDWk/jTTTbGDg0dIda9ABc02BQFpE9RDCJigD
vhQxGmy3n7qBgM2DWFmcyBdTovJXskQhCtUE8cyJ3/4+nzhubMKhfWKAuiADzlFZ7qBUWX8Vpul9
AbgKFx3k28qgBH2KuaBmrBTHQO+VddpCE2OZBleOdVbpKkyWdDNmHX42hr9UEbS6iZ0Gav6PBziR
2ziZ4yyMzOripvjVK7RX3f4BeJSeRlz24cOLp0uIwfzU3Nm4ycjdoyAT/NsBrQPb4/pkKotLTg5q
B3e6JqzjV4AkFBMz34djRp2+VN2wyXuIzv4vpgnsD+g5khhgLATSaRpVHCR0B1Rv13muYQ7aO6CK
LnxTltQB+mrbrn7mVyfw8cCrbpaXEJ7hlKsX3s/ULqS3H265LH5o82mzVxSKFELRjbA+hhauKBr2
p6D5giS2YdOjL5Dv6ayHSvjf+ELjmVOUiifCMcQ7dikmeyKHUV46Zdir+YPmYXIx8UEHgCFhXOBc
kRIv9R8Rfb/ewmScz22K7sHkNcHwkFvK31sMHoD8YTuRAbBfN3Q1HhL757Ity/oNovRnvEMD3Q6G
h9MW/m4R7fDA6Xe6BHSb+H8+bVuAywnjFGqYypxTnIowGz0ZYKl9isqW8JPdTRUsYROGITqTxefb
ypj1Pgak1kmKb2jeeBwMD1zec36GOsSMBYMGijKftAPwoqpPK7XioKSaRNRZmb/2RGe2Wx2fN3wX
+Ite9NjJJf5pncKJBRhtyFnf3IZGmRRtsR+SiQZjKj8Iio33+//BjuRy2ca6ZAzBtwvufZjE2pex
auiZuvmhQXoQHxRl0rxnvpIgLVZDsLl1Hau804ylZVhTmw1xGNTELUGalE3P/7Qz5lyZaFywedv9
uVH8uzuIAghhO99oQw+t0LCfHakxRE3NgjrpJnLkcizqSbBQoF0aEkNn56mq1DXMykkZk2Dqv9lF
Bzdzh19QXE27deXlUMNDsXJBXUNk18+3+SR3WT9kXomnC2yy+Gjm4/J51wqMrRKD5j8DH3v+DI0y
72ABKPzcX33m60zHcVa/7GKsp52FEOHeA6lSUuU6RawtNnITUwbofPe5K/XHwg87yXj71UbEG6xr
Fyj068jPVsoxws4MnnYWIx6OSUBphXP8f5PGP5iw4y+ETnAn7j4JIhCzAq8suSZz+1gyDaH9F2O+
v3uzddwJZzqH5yoEGvop9rYupGWi0mub+W6sOZHIH3rxbtF9UABxi5hzCkF40qZm9xnjeEO+B8iI
Lx/dxyYqllqaBnIl4Y36JhTAZrqo3ceacba9OYUNTr6Snn19wZaXYapvUzphQaKh7jc4ut4mzLm1
InYQt4kYqVeVPvyrisVb+gVG8Ts6gojBH7QGRPXl/yL6FUCNV4wWcmiM/zj9OXU7h3uIrezT6UtV
khVxlbnkh07vqFfuzIMjJVK2/NpWQ+krlRHR6R2odMex5OwMgV8ulio/gcDFAJAyrwozBQLu6hLj
xfKyQwL1OvSaT8mGECkRH5Qh4BtVr1lrMAgTBio52c4Ujx1j1gYT2kcjUc8FLyXRemNDffxE5iLj
Ir6MqIKv4XCsgNazc5Vm1azen9qK9vWBd1qoty9oGwaPLzqOtsDPfV+WPU+5WOz7WNtCw4arfEVX
3OIRY/Jcz+ksrW/oKtcwUN2ZM2T0u9JRpckZYH8kvUfPkQCRmO6vK+pynO62ynwrnTmscJNBNxVF
Gw/GmvAp94ntFrT6VMLQar8D/DSr0hcl65lLVwJobMH1IWBWGbw9mXg4iHc1hV132CDcUpIC2taY
fcTtC4ApTTv4jjMk89HHLJfAndILoJ3m/gbkbBaaEFx/zysJrnHs3HHvlJNVG5/bDaXwlQvCDIKb
6i/aHuKc0T7zoK2eYn9pvoX0JUt+ta8fZQnkQ0MIpoKTrGeFIIvoydSdR5UazmdVnvXc6Yu+YUJ6
0LLDMGGLEDje/6pD+XKi31LVq90rTcjVhB7zH2bpiz3ipiXA5MnH5x+bJ2z+rVowMmelrdHUNT59
+bAn2GxCp2NqPvLY5fAEAIZLUaz6Ewi2q59yRwrUoNhPePo1JVx79KPxd3hZu8AGd8QDqoewili3
WNTaNoHF8ZdhUYHG1CAFAdTl8/89S7zZyfuDqEcG8t4XLNT1oWF1YOSFY7Mr5K9CGCVsPZwod8Xy
IWC1iBfetevxHcNgSHzlio71wMDMDAQ5VGbTD+atSsr/9NEd5PLbWrbKO0PV5U89SGKc9q1KMntJ
W/ZsK77dbDC0obAMmvbw5hKUuWIPlpKyjli+oE0cgVzC/WY60ZhhnuP8k47hSSYMkGRxNDWvTzUz
aKfCUtGCKttccigKQzYUiU0ScKJFaf2Vip4cfzsQMQNnFfjNCS+6ZlXPY4Krc4uJbksQbA5oNnu7
yUWaGP8V/z+dpRYx/WEI5BXrgnXb1NF62Ltt9QolxS/GClm6LEx8390ce/MCNEFYfgR3SDCjYxQ8
GdjoQfIj2T5SRScoBcOCo4BjASJ7yAlkJvZxfU2Id/nxl9YaPqIot2Tipxvso6P2zbJrKLy5V//k
cJMAnrhdj8bjk2xzyGiKqWtoPEGPJwIYNA9qphaZ/bMmGQqwJ5QQEtxOZ77InrG3R1iJN3QhT5Yl
H7JDeOG1qVH8QjUAeE6FXN3JB7J9DL1yg4/C5YPbpPQHpC4VKnIlK6YWxJ080jASxtMrA39rVjWw
P+SfO1RviW4BRX702DEZFoszYjpJKh1mM+BVytN2KXygZH2R3ot5Ej2iAeOi+RmbNSxuTM+ra1Q6
m2Xo1u0WLE/tHRB7rpcpFoX6zbKQNw6qeUwXd1+Og1ZYru0Kt8/eDUZg+vvHbSmuN97kq3GQhHt0
2ruAtzFGt0oB9ka8swIsUlDGGfUWp7AjTIfmiGpWwQ2hCIrz1Rvw4eZKgFwiLCnnXVxF5p7i2Dl5
nzMH+te4zGGEtDAWDQar/nZ6bExxBn8yyQmQ0MzLA2RmIgSVdI57u/sa1qEmBGacgxl1D6+KLRO/
3o+Pp68dw2DV40WlbG7Skqp3Mhr9LTitp3HZpiSNdLz4n0xEzaeFmWIOFOVWc6a2XnFzrWTINywN
+aOAUTlfjfrxlBF5UZ9Yhe+O0DsRcKLXtNjifEVJOckFNG1AuE1/+xMzypB3r+hAxo724H2nKmQf
Pc36O8cEHj8wx5AAR7j5L3Do/e+uZ32ahLkycKECnH91n1IXhficNnN6BHmRe7jvGGHgRPh80X+8
oHjpPu4eNBu5tzvZNDejRRmaYHsQnBlQcC83grtwvc7RSXVTe0KeeMOUXiSZYOewt4nEYt7bqdsc
N5mgeJpTDDhgNXOx8CIA934PblGDKAYFSbjI3YLp0iUxr0ND2Iw5Xa5L6EWd4s8yXw7ZxRXJtlzQ
av6PJ+5TLw76K/JK0Avvas7NeC5V0nWjiNkloVaxtYZ3agYyQ7lHjZWRAne8I4hNJMgZZprtBpAH
4tXQooETNw+ZYk5J5/cwJsfOZYBZWKwzTbNQZeP1T4tE/ZqYlmpG70F0RUGz15xquA4AKpTbGYos
2x5V/jg1lwYhcauATY01rkHO9tabCq8wbTDvSVS3ZzFVZMlUweKpJmYChCK8I3Lv8xe0VMGeNblq
SehEPtoF4efFfuto8YSbmZatK8npHE1F27ppzz7MztaA5/ZpQNkZVxTG+Vo5Xz1OkNkeV5hz9fwI
Mh/iWxRxIZckP2tSkxHQuWYKCNdI3VE1JwvewYVem2rJxr3dv+WenK78byE6QIXk3OVW+ZC4r7O3
SYJ8tj5M6v5WpUjDp4vMZZJK4DvgsAuQn2a0Lu7K4JxW8Mn5Ni2c2EUG6sl+uII26y4H3DGRE/KR
d729Gy40VMPQtmnzijVCpxKnBAGTTb3Jm7T0vJf94WP9mHINacK0HWe7aNNdsYUHBfSR4Xh+nuqs
l3/gpcsptHxNS8UwmjoWnLJ/v5cIeyFpv94Gxfm8iQHAzSswgaBL52phbuUuAzm3UVeTgtlT2NCK
2JVSFqscs7u0ZTO1CPXi6+J9T/BTBBIMnoaHgiZE3RdX7CMsMoUXl5SGo7WrntwERJq7elbI/UmA
aApKlipc9ghhXw/d7Jbg7sBSEHPDzGAxt99iq6Ui2BdV1CSS5GiFzWUtgZKG86EJQ06mca1ajTvH
BNZVntPIzMl05hAworyiNkpIl189CvPzxTMmEv2jNOPsU7fln4tPamtVifULmSFe69lrYXZoBYZL
BMZbX5oWVRTyjtKugOKghq+usNRfPuC0dePA6HHTc2X4+EAUIDz2WRnrrMKjKGc8iATBa2LvhXl0
Ifu68ow0Ve/5a0GMf6wCt/+2+3qmxvyorSj4+2Rsf8eT/EUpEa8jQM2dRZylRhvs00aeCmI0kNFF
VgSLydbBIoJRK4kYtXZKjc507oPdwHD08Ag6exBWx7Je/C9bTuSdAtrfAATCHZFp8uTdCjMaW/8c
1rQV9TetbtPqyKSzxaA6INchb9Kx8Lqq2LXxTXS6u9iU4+iPJIJi6UKpoS247iejvIjeBj/GMjDY
eaEPHoKMW6BaHRIiy1+7R20E+QbGru0vXlDA3Ic44tNPAS7D6ewdY2cBsfynA38e4Hn+n23EQ8Rs
ksD5HOJZ6KN83csnjJq76fACZQHrVRv73YBtAQkCNbw9YaRCFsAWzpKQnKNlSa7+DK2SNy4Ytkfh
V9w9zcmBwKR1rtg/dCxRhK2yMRYl/QjbBQu6SlNa3PckYAmKlLSCxIAhZl04HVOJ8dXQPcjVafFh
+/Hdf4fT1Gwjor6EE1gTMvj5tEE6ZB4g7fb9mBGfF1KJR1st3NpMDCqJe2QTBN4Wzzd6GZeRxR6B
0Gh4Og0ss7dzIhMbHuRcSWZ9MMdMu+n80HYQEDeXQ9HMro9dzwhtuL6YM+90WN+Q3O7n3OjVxZnE
yBLVneR3FVehLaNP8QokYBgqxrKPqOtdOIVlnvOZ9ILGyoUnrGsR0lcuATfC0+i0ezaveEGy0Awi
TGIqnoXGpO4oHByVmPQBH+ZCgaZofy2arMLVDFozQ6OsmekYp3tYZokqfVYp4AMuWYSv14hffgP6
5CkHC7WTo6xNQN1tBCxVHRngt5Hv4P8H57i7rOiDCkOqn7tpjPrqU/eh7OygRTsxtwg1MvhdTjOp
BZr4aQury+AZPiZw3mFy2ojB6dDt9Zp3VGOpDffvhhLJ/rTNyIJTTgQ2wMjO5u67FBAxfDFZIR48
79uDnx+7ep+IxSoyCsakxLwYwFjkneJskueps3GIyP/pyqvShApRS+3vzOMXHcMDG/f2S5SNg5hh
VN/L79SHsedqSFTgR6tmzVcerL7UsR1QBSaIvn3v5xOqCPyFted/VJ2O57V9QL64XF5G/NHLoxww
MRzJWKKYWXiqT2Jk7rMJu8LROab1PJ9P/UgcJbhGPUnsFq64tY7ctTAFbU1EQa/uIYzxCbvRkDT5
iUGwDRSI5QAo3YyFmmLkNjwJN3/GK/99GHIQRZl+gQaa8yE5918r6nwlexqUqhoR8/h3g1BZVyOS
C4NXIr67teREWCVqwYwmsPfdgjh7DaFTBDPwj+4rhHeSOZzpdUOBZXCYTo/HtiBR/8XbQjX8Iilz
U2x1u2uSjXZBtw8aGfgBjApw6gIxCTq6uWpZJJ7kBAnsW8JEcKAdgJTKdM5c5hoXc4g8Mgyrm2U7
VnBNuRsVCkFKE3LuqvdskINcOdRuBZhmLoDUxdwS8H153j8HSYAfX6H2pZZi0whQQv9dSkdKbgRx
+tux3+oohmJ6bQFLaC6t7vMDOdTHtk8oQcRwd8PxpwqGIhSPaFkmUoLl5R1e5h9rSDoV/tVBBk5t
P4hm/l3vk0VpHjk8wxCqgzwqXORq1TBI5wY0ZwiMiofyPHFDO7tNcol64Wo8+3+6U/KxMatkIkC8
MiJu70t9yQLFxNy9t7noXsFUC38Oa9eGobckcA/QsQk0+eCr23wXzVprMXVT+JG626zsj5M93lxw
c2E64SHwxA6hq0f1/fkcdqa916MPrupowaBOeRTtdeaLoI3zUxH1GoPEEJKEAF0k+h215RpwcwF+
s1dmMpbGbrHAihc57FHtOeDcGB7mcvGg4uXd6A0oRwHnESELnqbFNwR2liZSZ9jrABluyY9socVy
CPUUVps1LU35chaQLXFkn8f1UeRvdVbvInSk1qd52XEQUpSe4DHa+qLW5MTq40XTF+iCt5j5IhcI
ZI8AcyIh9HksojjbQy1twdoYva+ZTIvPQxkJw968b3O8y/JvRYldIIEnstpXhm3nzDfYu6JK//we
ZQN2XjnTg4i47k52uBvannLIIm+37ZxxFXJ3nm93M4LzSWg8DxNobIYYdOthARcuZesbCssaY75/
FH/9JnbMGajbZwKbXHm4IyCIU2AxSsrla+nIpv686PxqIPnFbm9vBwhvVY0XAskKSMBmonD16Inf
hB8mfkLjYVvK+Iu8TJRnanpphDVd8YqYle9zg4g7YzCSt3tj1SDP2v90aWuvrHrGrlae9S1T80GF
VAt3sBokCWNR4gOIKgTtB5YfrgUvAvkg/LB+aRIQ7eUPK6IeKfOZQLByqM8OZKJ67hO0NhgD0mE2
iduQAQ/qs9o0AzlaSxt/aXDE90PlShqtaxmtnuFzjp2H1Di4IgOl5KamIS1SsCn8AR8picHEV2e3
oZ6II+MnbFaCEgxJL8+8V+qvUMiCGnJ/Jti27PXkBsBGXa7QsTGMKixnaRTAvVWLI9Aqo359Z8gZ
/os5PHAcOiexCuogYxtwsC7743dtYSTICAFeqNaQMwwu5CcZCu6ZnpLQdWEp+uihKN4TS4H7zox4
QvN9nk3ohOxnYlIv15wG6kUH81F3whusSyOJPVzVVPQGF0L4Y4jDvLDGK10Y0W/t2U784fu/nx0Y
LazpXUB6MbnDbressFfxtUCP9ykofAiE9UboD+CCUOu4+tQnGx+golQyO61dqo81sAcuysCnh1iw
+aBp0dE5W8B12j/yaVAxy43k4hl1Nv9dSsAAitj4UwVk8KUw9x6XSCk+fPirVUvMSh0qFHRgZzy+
em3AhhyLksXpwgdlkUB1e/iKBknHOfBHVGaDEpgX+CfArlqpYYBViwLswtoGzyF1sFswPf9HJJLG
VcW8imnTABZxdChRsD21+klemF/7ThDcRwBwwBa/6djlLe79ROty2zWBbQqwUAm+CjQZPjLe1TxE
qAPrhOIuPQR0EZxa4l+xe4gXKu8PwZcWm5olA75umVmkLWRKThFnGsIgzvP1dwjKx42LJCKOYfmS
RZ7Tc5w9eN5I2nbquVxiDvMydG7xWeL2zzlAuEkx+j0RDsQY8kaefkeT+XODsexNtG7Tk52SwK6t
VbjU4oA6gBu4Q3wz/D0jzWzlv1Cp89uiCQ7C2Q23Ebm5OGuKO/SEfQhBRbvBrZQzGuTbB1409J4X
SJnNYQ9oBVU/7tK/SQxyoHaDorE/mOWDz6BynE2No5QqXqcSzSdYrjWKuqhrb0CTWgKmWiZLHtXD
yP1QhC3VoGVukIcJrOnStC5+3slPtb2hEkuz2+Xlk4LUSM1gNKhwWbT3kODbDc/aO5nsbDkh+S+1
d/2Z+Ku/dMFuGWMaFyRXpZJUz6bEVkqjITZGQuHM+be8VKLKWDlPuu1O43Pj9aTUBWTNKfjrNLRm
iJD7N/eEZ26r4v+Y/0+n3SDL5IwC400ZE/r4zMR4KSbw4Cd5AbaFSN4uZQA1SdzPvcok2tE5nFce
slUCODr5A2AAHuRdf4ZX1AgSOXt/0nMZCd4KUK7IVYFdOs/JmInnkmDwcmS1Y6FIZMGcyR6A+QQR
cjPQZQ9X8xg8uNx9IiQKVaeA551YA+LLPAWgxodHuNDYlA3ZQasy12yb7xCKXPHjyQoouR1nAIeu
KW9Thk1A/phXEf0PsGhL99P0lcQIyQ5okHdcDZCxMfTzgb6HHiDOmzV/lrvMMcLeGU7qXZIqGPHb
4O71RDtLS0SexvZSxPM1XfPT1zl9l/jhiCA72hNeOOXEYDwNr4rOByZYFsndXcid7KUTLYlvWbJt
UPF3OCjl9kt7BPht5RsUc5QPdRCI/7Uh2lqgGcJHryn+LzI9m/qnoSPuQqqXCL5O9VQ3EQqTTEzY
0OFXYd7RBuKEETUx8CEHQStKRhlD9HLCFw9U3ZyQp+raXbOTDM5qcI940g12qc91jDklHuqGxHjP
7K5rSEmY+yJ3jLJcfLSGv/BwxXPsYkSu029Cxtz8xf4QnJ+RRMI2J2yOTurkNgmiWChMJqsykPeo
N2PO99ko4iMAoHAZfc1kR0+OdlydkacY9fke6RW3B7KyE+RcDUjAULYmmfrIV06E/WgKendrgNzQ
C617/hffcRl1d/d1Pr+UuAxyA6bsMYxPDxr4a2KGhaLIUPeZNnMincApQXFZn06g6iS3ixbq4bh/
edNVF85S+ZlraH8JStQNZAVl6yrbOl00uprXoNEvKEQ+ZYlClF3MN99JdCPhsG8oVzP0gX97Z5Vy
KkwpVMxhLN/zBec5h7WEH2cdTMvNExJnnrG2rN5nOKy16VLaDCeSne3FQP2c1m0iB/VlmyZqrXV1
AF/2ESsDR+IbGAWVkEs3Tai0bwqrI3j6Y05dfq+a18n+E7Lvh793iVa2OueA5oy81WIypuiCEBUw
AIkE/Rmgl+ufTNmW+ObWxOHj39HGtQOrPzZtoAJeDe70n+n6eO4FnXz9smsSysQzKTQdphAg0x92
Pm3sL12g1dv99GbJtYqJXfYbe4tRSRZUrNOYa8ST9CjDkolF5ppu3YjzxKAqwmGfHgh2gUovxnOn
kEtHD3shzx4Kb4I5CWjQCu9EbgLytiF1ugzfXuwFXUp1iqCtmdTDsKRVsDDSN8hE6fQgHKctsxHU
maD7JgqVDALFv31+HrC7S6qK01OgaTbtvVRjGjx+Q+b2Pwul1VYjKvmLrvvU2Zmdaj0fDdB1KtlU
wvGqm6YfcIHqhwqhKpV0Ul7TjZUKFCR1lrzG0uh5Ts0qYWjk/jMR+XBZXIPz/9Gslj7CAV+roofK
dwiOT8qHC0HAfghEt7yJQAdV86tsZaxClFSH2wPBgZwtQX/R+GqYQeR8zFbFXNTDvbz6inHhgjEi
jVwac0vXVFU9JIb5tznewHsY+4ZiXteSre3VKXCmpQWsMnuJBBiWX/l9+Q1CwyASxF7onPuHeAgu
usfDQEQJjuRzEIXTD1k4xOyDy/uJzJb3kA4ISFzh+VuyzbHnd7z5BbRrLoxbedXNYRTK6EHyRm12
H3JDKZ6XSgii5wH8BnoTTH0D0ooPtRZDzf81xn396I5LE8IMC5CqB6KmgnR/Gj+BtbZWyUOuRdnX
0X67/Jgv1QBRD9/SU+IfiDo9WlPk2dylEBaT/HlncndnFiJbSJbmdfyq3InvrCKJSIUiFb71muzO
DI5/rhlWTp//7kqmtqUs20FwTZ5gtTqeR+UOvWh6bvtfhjzmIsfxpHOhTjz47pNWQZhlhEuR8zCR
h0OvsHn4b09E2LkguJQZ9OtQbPB2zTYtckdHqkd8cAP25bC5XpAQgc1lmq4LjVyCfMs4+A03uOR6
+aaRFNbRc6jnzFH3SCuSgfPmFxNyFn9PQVRo8TQIQIC2BUC/3Wh9cCvuxHQY8RqUfi3WBvpZbXyp
TsPwFBu+gUS+33ju6bhgmKAmKvz15gT+2rrQc9uu250nyDmEK/ttEh87UbX4CjneDvBh6TO+WUC0
uo6jqJYPEVNKutsSkFERAeZJhyoGZzyxe+Wo/xEvh/g99foDXWmLg4wixSV14nuTXDcHTbVolYJm
IFe6WL6YIqKNJ9uC6dmDPAZ2KZoK+NlxVyng5XWuWpKemdWpuuVXXdTvpU5BbzZlg1Y7GxxxUR0B
xx1Au6U/A8VPciKsOTj5EGSIKHK8mEri80TfLXLhVk01tAkb8ED4euiKSfK+kIsCdCA34m0eInwc
GC/WRmA8VL7aAsB2kHjtWGZjeo059q4J3Y83P8zDAQ90XOaiOIJQIKuPHcymgeyxrlOntf+O+rH/
5aFvuxXiuLh/PQ05vf9xT7xeE9Ere0WKNbyJ80xs1OBWT6n9SULthBEPn+35MEq/fXb6sNbQYKb/
rDLzCXVv8bSO540Rqu4879jhz8jO4ox1pcGAPD03rgwFup18Jofok8fUYidVObBD/bdsMZ9+MRqo
50Y26gniMkrbCQmHtn9X4KFY3cX4GnHuM1VgUfq6knyYmA7JeHv+Y6YBUvBfghitSlq+qdzoOPIT
j0/WPXQv3v2LNyM6U3rO25LjCE2i36uRYpfdsNUg/PdaeUr7BijPvemJh+Iib4AFyCt2eGLj8bqr
n0RBIQD7ocXfXfYXaxGXjgCPkaQcG0+DlYmz79xtPZn+xqiKPLF8lFFqdbEi/oSmjUr7WBADgI6X
oBdV61j+8WSsxHiY2vfEDylr0dh3U4vPEBqSE6ASBtmPNCBJQbRMMobDLaCH7R+5sSN7X3W8LouW
U/32wJ2e8FB9V/RTaKdSWpAM4JPvI81ksxPtC2sGORreWGFjgeKj6ujTazL5V5JnNChIqVK0F5K1
8gDLPYh7RZ1x/d0AYDSKPKxF6Nxci1MwnsiUGmDx4JwiL5Bq7hRPwzvzfPTXyL+xiazzBXblGHiy
/TeB9lx6DHJNJ89w51XQC/SOBxWJ7zrdzBGcwE5gBqa9+oPRlXMFPJC+X4RMtBkRFgq3bzP0uxhc
HJeFPqSqrjPjLdBQ0t02CCYOyx73eWj8kM9Mb5fnFLwSX4YVGKXODMueNFiR2N7YkzV/ShMw75ib
86AE7NEwZ4gt4sA3UURhUFYdwq5suN3Ha6qn4tozzoG0PurOSFarYyJtukFQhrj6E52TCA/Z2ejE
IPCWvWRVmbf7RYc/xapEz4aWlpxyU1ZpXHbLi/U85Hfm3ogcla8pMUipSWDxyABDnLl9eJ32ci64
VQAEOKcXP/IaC4vV7m+5mPeNSd63eXiq0EQwcE6FXAQC3XnxSkZOutZdtil3jRZeHUwfldGocFc8
5ug0rHsbVvnhptu5F0/jTDP+OrBVKdBSkjjz1T9QQmuf3qLuzL4EBCJPnkM6oXB82HNDy9Vw2OIF
icuiMRecohA/vaekUmlZUgfBb6tG8XXresvX2rU1GfsZUmcAHltZ79Qope90edWOahtmnolgqaMd
/ShahLqtDRaaKKYbT6v6cbPEeroKPXE6miHc4RiVa2n2g5NkQpUrXi9/4fRv1SdLH0q0iTsZ6JT9
ntPc5aauBRkiwxeouBs5KmaKi44F2GsQ3VvzmJ3LcnK7iSckxGc4ALRmNWQx572LnF/UcF5usYDz
eg5De7vnT50+mVyhhLav41N53bn02TV+icdUB+A/mgmE80VSVe1PuJTsz7Rx8STOXHSvmAylkQXl
CyS0ql67py63PdXXjliFe3ypTZaZzA++ZAuvGqdxFwyKwW06hk1DcAFyqDXckdpKPFrJCs50BOD9
EI7V/kjjySsd4z8ZQMdDGCs62aIsZHiIL6tLb9Tcpy33ZZSB6ePJJNY7cfek0QMmZ9ZRf/FPX/yc
89M0l93cOYCsjFDQmBhedgH9+9EbxcewMoa/eXXM0OngOFDInEN80DvAen/zfKOjglMwcXP4ZlcB
eGh7z3WguDB5ZO+U8EpyN2CATv/9RIjm4U9+daM6vR8yzPrXitWG26armsNpmR1ZkMxq83oRaUY9
3BAA/LI9AFuFsy4MaJJ5SnDFmrA9s7e7jIaXUYTPXlejIHZklY7UCI+Qiz2DxGolqFe+Tc6fxvSB
P8sFCX09BHGYBVwYnxhadkRSuNgQOuWw6QUa3IHepPTBYWhP4QP6aEBsYZA9ePVyDNuxkqmGXTSy
uQ6dv+Eqe8XP7P5+YdrNDziK/7RRYN6N6yJCmSeo2pj8tsq2aY8UHFQKW7gsC4BxiNV9pKq6Ob+V
inw9Q97czy8IdjuWRcWWuJKfJTtb6Z3rYKb0r5udQy6il/OZDG4bLz2/U0CgrzBRftRfAPVqkgNV
POAJr0qIjKrY0EMJuftUqhGbjx3FZ3B7LLa+/ur/N165YcmCk7zBzyzwImDZIsGMDxSwPmC4aZVW
Q/nLJhVt0CBajRFBuOgCMxX6BkAsT13w70rF4jnIaXVShaPPJRamqSA9d1z1FN/Itv8E6fk72gWJ
FIKJ7Pik185HQ+Ry+tQO24iOOp2FOzmGlfHjn16f5+aqTMoM9GfGgYzN4nTiR+ciV+PofKHqLKpf
oiFIvyuYAX+Q+CCmQbjZ51nz5zMehq8QyqYNx//+MNC5cgDPS8mafxB4V0HwGudevpQ+2DBmXeSs
0xRbcUxr9eO3kNJwkuNZpPF91Zw+CtLBPEKnoS0QGYQcj6XeKiHdP7D8T1rCc1jvo7xiBv1zU933
VNFTOsevsVqlNmBabQHHO+H1yj0vlK2s0jenQ3HhZqu8uhFl7vVodeF17HswfMIiuU7GSsPcFJJR
ETKqNBnMD5y+vYnAI3ozrtJVGB2QUFRHUQXBTpyTIg8nVb4ANfG9KRDY0vzPhr20TYzgOrxYn0G+
DFl00MvwlWnFP2BsEWzymC6+nRBw3+KvATyj3auLpbuHQmUiENoiZElty4zfIgOnXt8JvjMrshBI
eMseo8uOmPwNgzwJrGZcmrYhZ85IMwwG+JXJiPkThlRblh8gVPfyZAmoZ2hwE5P5Q0P0AkgRuzCm
h1c8bNDP9xOaOofLrMs9oRCK4jRwT1JeEm+puFO3gY+dBjZRaeLpyceqifP1YoCzFILVT1fDhVxj
+K7HLg2mJIyq9PiRhjqZCTq8mo0zTdsY4ICg41VgwyzX48NgheR+FQAUgE8RTtPbPtQUyASdx8FV
hpWThmzyJrhK5hXa2N+i453rzxxBbneQlD7sRVf2bP79XuHHMsAf/VuMPKLXJEIGPnnvpCKBl3kC
HatXoDZXNzVHt/GLgmJKZpMbHpPfdWgY+EMmMgcxZZPUBo8F23Pr/IDK2Owj0U7N+HaxJPwpqOPG
b6eywkOOLKn6bFM3NgnjE0CfBAcRFrGd/zfl450gO0h9BuHaFpjSjQ34AYPfJ3dCP9NEZaWHiCck
u5rxv46pde+c+lYwbkxZC6LllbTQ01CPXO+nYadsVy653+yTKk35L0j8jL47wv6jmnRQ6euN3J3k
4dGUVNZINxD9aR0qdfMv9Bc1mqgYWgUY/iiA+893vIbRLzqFvypqvstPgZ/IS7Y8P1EKtkwO52mM
etSH/iAoYEs0a4/3fUOa1MN71e0fMRuceX3EKaY7jjagJqlmCO/nnGZM3ppD0sA6NBuXF9pfYxac
bDGnFb+MKDUcF90xfk9sagm+jukSISw3+f1Viu6AB819DD4h3weH0tu35a0ERg8P3odqhOi81CKd
aPD1HHovHbfnayO4xEn8kNo4yygEcO1R+le+9JWbu8q8lqR8a7F1f+LXTsLByJnxfnrKXAYbn7zU
TnwcqnS05vfnDUQmGwWKROG4YA01zQd+l0U9HAoOvknUS970r7Kl5FyMG7FZ47zoME0FjfkACixc
BsjTYwQIqrz/aSqsrHadXLXCMxIT3VJqUKVQ3m7C1kUy74gwV3Sb7AeYUFUYPO0SVnUqGHCc+YRS
ElnCymBU7/vjy6aVT1BrmR7SUOxC2iCw55s1F+x+rhdk51AXm71avxVDg60yzSkt9eZ3V0xSpsGq
WQp/GdEsPS+sPZK7VVOQdvHNZuWvIEJ+JkSVCTRaD00H4rNdUaggjFTzqjeNjlJDg2m2HqKzlLLc
cdJZv1cFXBPV/kVut6EVEF9QrjW6HBk9mFgTwuxBuEu5Kh4F2RkfJzSzX4ReokMx4kYLLQTAUT84
bHnFXa7kekIj48RM3JN0n0AMsq7j2+vUP4ZS3sbtQPjVLgwxp85vV/OIqCiWdnuhP89V9ZJQrbsv
kCYWWHTKQC7q92WW4+xS+heJik0w4cutrVlRqF5Ry5c5q13n3LDj/lWUgWL/Kr5LjTt7GCOc06Kw
mqmFeBjrWCJkrYOKKCnQr2QAI6Ginm+fby1sTF9mj98OjePNeKB326eoEBxew8GaG8gA/S83ihm8
DpV7vk8mnW40sYMiF5UFylvNay6Bf9+Bt6LYcUGdcPjtKtjs8LsMN0Wq0gsHXpXBi4/If0TkYHcY
WMZCmviQwjnO5Sv2x6LbHVgBftttwjB67YESaLBn1xYLTX5RyIh8w1vFeUobcgfrJ7bjXX1ZSGqe
8DoPmvMEKs9zDC9+3mTZmTYJ1wliMvraXm7SYfpdU+L3zIp2eZ66u6CP8R3aFpyybP/GjmkXdZtb
Mmubm0GIkZKJXuBNujgc6OcCZtMYUA7/5KUbCZlRzX3tPEd1wrpNE35PNyKZ4GaVeV9FHgwYAiBk
3giN9kdBM5XN9/eckcWmhPjI2+mpJPDAgzVii2dIlnuVCIzHzZBUuaibn9Wbsi6rA9lKZq+eYDMz
sATjNjo/G/mOwaIkXM3LdfBGmPnenLQ70DAL4S7FbL28e4r9WGgImZdYRoI/X98b+g4UQ2PcLyyT
7tl4yjQZMXgryD9GGmrEznsYQQVqY4Ts5mmIK2jKSUqXHlYX5KWwKbUj65C5GV+vCtcCzpuy/0Ju
JB+GoWsEAJmT3rjvPB4zosSm4WmjjDnkApZ30/u3nP8EdFPthROqCoCJfWIu0/RYgzVdQA02WD12
Z2M+p0rN3zUB2FvhcyLb6OgrvQAl444rANqV7hUbMjcOVtXUREV2WOtwl1wJmKL0t4CttZe/hN5d
pw9ezbzhU7V4eTG50pkQK0ZnmjDZMBnaVxeHtweKMRY65KdE6OXIz9BhMiu/3dXKsiIhXkiqaafm
LIvO5Rrm2BgVFw/27+XagfYQhaaamF7+Zp2nMLnhXksJAVAQzsX7Ga7pARUNbe7GT05yeeEeDfPc
mLxr03pC1qe4jbElZ4fS+bIg+4DZDK/PAnnmwlQ8t0sqW1YnEgeAkx+/GcNuZAC7NizxgcQAQ0e5
+dxK5U6T0fLkJiYx8v4prGDFAk581iQLlkjvMNxKaUrQ34iL13vuE+b8z44rCVGFDrJursL3xzUw
AmQglAc8amm3zxWJFyvmOSowXJ365IZg0peamlKxmUBVTkZDvGk4yHo9b1bT7QmW6JmpiuPX/eLs
MxOalp0/9KngDeCrA4I8Pp3c+MHIp/nV6gURTrZ8zZwUFmmjM6fPOym2RI0DCMzCdQs2fJXDbgxU
0H17evcZLy89nsF9ogA5tDL5PwwM9Z39MIZiqpMdX/yXOKiHaoeLxS8fPuVGjRkMj9xZgobs+IY6
HzbLygA/F5+KeIr8UV+2OlzJb4knDZYl4hLzSukV/XXObxt/vFdd4jU7Gi/V+blW1L4yxXiRhHv0
zMny5TTPU0JtgLWVW3dITqhfpNCrFt3Z5tBgyyLYQ5GTyeijbl0u8ZjTYblHw8JUALioO8aSTSFG
UZS9FoNZCIq37C3KhxTulKqQ5qcmILp6+gi4LYqRAqqw7c+7Sq4NR4a9fXVTADaTYBGf5O4GQhle
srDKlh31NetoVZFfRcLmRf5gJ2BRDi3BJfqL3lAcl2SZvnJzp2uTX8nc/RBGL8WbeAVdTAN8HMPt
EgkGJsKaUkPEHqn93UIHao8ScaIhl1Rd5hhg4T2cBsqQ8MBYSss5AFMZo5zOeIslEVqaH8Jr4/8G
6+kRIUAiVIpD7e63X078RvpyaVgtLVT8Ms83ynRDV2Qoh7V7z4kAT5KAO3JXYI3ScBf/cX9MQdCI
7BAl2oQtOcy+l7OMPbIBPmz2kqzHJJJp8HUdMxiSxzizngidtu1fCft0B/0vPgOL2Br405v1ofDg
3cPd7Cq7uCrUYyzB/cfL585Iby3An2HbTWwW9VTpilB43v7kcHdx3CfQaXkq9racm+N2Rd4pODJs
zONN1lVMcvGo+9kZJaTU9WbP9uf2WsF6NGDKW7wFz6T+6UhUj8nEHo9Y60KUk2dxgPT27MlMndIO
ssTVA7hYfY8QtRbwwKlPM1xhn8UuYi9js+e0EUf/tXWBHTtajUoibgl3lnvw+R6vXJyJLmK5eCFR
eTsEJFpi19SlugFTIo8awmH2zUOkzIONeNblr2HTMLM2zk8lVrc2wcpgBguQDfL5tO8TIqO1iJQc
+E9JDq0SdQvV3r5LalBo66g4GYY7U8H/qmvsE5a2CK9tGNl2k4FXaoCTcBugx5m2Nx22jRRIWTNM
kCHjBrWZzCvHIh+jxALIICIHfDbwHIzwUfdNcZf1DtKXX1D7Qo5pGeZ53NpV+MVm0lUGFE11uEO7
OTh2DpswcQUBaWJTnc4TDpol0vGxdOwGQc5rRmWFnyHTFDsuvIjeglNDCxCcaDWYkkiAAxD/hzCo
pZmuf59HPIQKOaVC/P5vxH8qUs6AOWpsmFW5Iu3XRPObJ5a3UhEV4FLdm7s/AdwGnGxxUy1Wf8R0
rZ46mffLEMdudNbphOoKxPlhBOo9T7Sskp4b4BYsO5vJvCChkBGEJsiy5u2qv5o9b6UkuTxQDPWf
iaBB2tZAmxf5AiYI7VAHbDcMXit2BIDwqgepXR1V/bwgYXcGVBqshHqwSKCRtnUpDK/7DrIVJYSD
2reoph6Cx8wcMhCy29Dbld0vhdYx9mwZMDiyjlD/CH755DcFQCZUWp34KF3GOXJlA9FGSkSCa8Rd
tcufnvarpvZGETGr7Z5Uf0AagZ+mLFnX1yUMLd3ObQDAWJuGpz5RG8SnAqAG8L9tCiADifD0vayN
yFOxOM7ko2eSEMoSv1cF4HjEknZf/ZER+qIrsvmvSVACBy/8xg5tKOee7bS7UFKHlJ0CDJkBRhbw
rqvbxhCbkN2Z8Axiu+RuaHRa5wPTycvtWjK0K2W/q1oDFp4yS3HEDJBYMcaoQjuU6cDpJNH1S8In
99WPmzaZvcBAOouxpt7mSus3QR8nNlcEOpwiibUpD8S+OZSX2szZQicdvi4mUE04WkiEpsPpNx75
IHO7HwJB8UVnNPMY8LJEuYpl4n9QkNbH6Zp3nIE3eJEZmFXIBQBjEsoTnhKjeAmf0dRVdOu4TOuq
OGBYG80Xrew4Ftz2RzP8pjKj2WoAO+dhaVZ2y9UxwmVMO/H8lPtvTAoKrc3WY+0cDrc5CVEXRqQQ
ashfgW1TnRNLKBukFj/bdpDt41JtCrrlSzzhoF0p4zTcMBO7tw/9lj9u0e9uSupWM6qVC7l2HvKB
j7B2PYCg3hJLn3TN8rrFgxO//8AG4nUA+Oh5tnBLmUpn7HSAvsHmnSXyO1CpvD/qXde7TCJmJUpV
Yfr+EgIy4TIm3OKbYf2yVl7EYw5WYVCM9Dx8ZHNFZ1OShcgo3XH5udmXP/3r5GozvP475ZLp6djZ
VIzXW4hszOkKxTqPcIkDBhh4yKPDGZGWPKwEK9gnOD0IJJpVVsDr+TRb5zjD6qfVxNbTif1fAccc
8Sh5ApviFIWdM6E5fZkayzkNnBwzCB22qyHp7XT54NKMsxLKVYRqDQ5N9pa4ZW4eaTC+yb9YkAi6
fslZfQFVUVPAeLpLN25FFM194/PxQ4cpUxHN0SQcrsUvcLORL9F76YA+ey0O3DSNoWXsNnaAub9C
dRJyPhj8qy1yCryL9gfU4mXGrw2LmiBLdY7YjhRneRkMb0w8Mt5EUCjrLRzRrPdWo3OBb5J+VEi6
VFqT53pVVETln3XXgFnQDBekUQXPpw0bq/p7YmzkA2PDGwQxg9ltBsv+/kZnScpiIOkrKYYiw8bz
jRomWnU+OXWfFGpRerF18p/1X6Z+0h8T4prbifxxCIUrmV5us5v9cc7rnMZjPx6TC/EuM0T3RYyF
2ezOeu9LYEchbt0m5m8mqBQj1m5GQ/uPp/oQtqOLjNmR0Z5sKm7ysDcclwme00Blg2hjZ+lQPjix
7gfmycU9jgV0UmjXn6SMf7FFVvTBmGYLh4qdaNk9sgIUOaO5Mmf0jXI2Z800d8FyJ4hVJ+oxxgx0
urcxgaasK62me1WwadVAtRn4inet7h0wsHj0H9v9dIdFDjqC8P1mXzxDasFjpGZXCOcyRuDKGJYh
DS2yF4NAtDvo0YfYL+Y2Et4bACjh/qP0TbJ7SGH5ocv0lENjSlQ9zhcNzj0McffLaOTeEEiyFpsT
FncyorbhuKaHdZ/L6StvMQnRTDhkV9e+PSQ6TupQk9YVRIpSO7yPHhRPnZL90UzfJgyDmuHPD4lT
L+fpn5dw08Ub8nYs9NGKVvVAP+eqqMKnCualog8iAx6xebhrzvaQaYaXhNjZXoC3j/eph0gMj1oX
WkCNylaGYkG/NBYGVaSvdcc/99VWP9MBJqshwrNMLCee9i+ydk7mWikyUvrQytD9w31OIiXk57y9
4Q2HWf7aSs/FUKSb64PzlU2vEr0aGKWzXuo18O5BF28Fz8H0zHF0NbB4etcoeDoSNLl9ZC0sYbVF
JPbr5CFa9HYg2uEka93c1veGHfktXoR6tqxzYHj3v8sRQkAl54MiLfr3KiE2B0QnrFOTc+Wsv7Xa
TGYLh6kNjbmRLDZ8FodIll/h+VLOfs+uOHvvGgj3tAjKLZ1weEyuDKvr+6PbUVRKKRB2H2TveNKc
gDFTZ9/VVtNnEJ/HWv+IxMclZjdJeNJHDdyUeqUaoMZWH57WcjJ4Uasjf7eYSRmTTcvgVJiOWHfS
JlG8qhW43CdmMLHLi7/aK39kdaZlM+quYMR94XTYLbvWUsp+3PV03mznao0QsUJkq9VAR8V0qvbV
j+3tpdZjPn2pidZq35q7x7ScJVUTjGx/BN4Jzbr5NL/VY42rg9lFbYlQMeOCEebK3F9VfBRxNV2I
oXxWt31CdtgP/PRE4lgYKglGIE//qXQigDjheoN4AsDqF3Jnn6uX96FLYJ5fLEnlifZnVkcaGe14
ltUbHQBUuAaw37TSgcU8fHCQOro2wpxM06EhSHD5eHIWxkPVVtDgk+7PQVntH30DY00zBVZeUDDU
S35ZtYETqLjRrmRp+4fAd/QK1W9ogVCLIfrRyoGvGaUba28EiTgIhdIQZhmnjGYg8dbAab27J3/I
+nWGNeN2k+DpLNUHeSTBoXZofpnmncm98ksaVrB3HNcIqsm5q3mY0zRi2/lT0dWkERoS9vHK0dkr
saaA+HAtAGmf3ftvTYvJvc7LgWhx0pV7Dt7pz+oZn0Gd+/nD+WK9fSsWgdLkHZk7QA86USbu2a8a
3jj5pMOfdj0OpsxzsDuB55RqcWYN/wjqyG1qf9GpGSymxOzUnq72H114bJfjUbYIHkQoEYaRv17Q
PGoA/iWRYQ20I6Y/fqCYxvHsLN3rcWDj2KTBjnylqCtTxcPP73ALQy58lVaJXCIFa61utsw9Kp4d
WNDMzs9b81KvmfCbg9zCF7QGr02AYNTqistZXPFmxzNbGkSQoHcojfKedaEJDtYkFqCeo7E+UnKt
OMVsygNTprLNUHIc7YRIOVi5K0MzzWWiLkQ3OeLfuyG3XJhOGy9Zxx7j61KrljiyUHApBEMAsVUK
WMfHE7uAV6HIF4ZlK/2yM36uOwS2aMJCDS4jj3w9jVWwJWCjVeSkrgYWXx8876hDp/65c+9dqGHu
EghFgmNDokw3DS6vdrG15Vx7F0Kyw6Ex/Ip+2XdNTyvn6tXceUIMNbIMZ/Ez1UqzVSQmVYn3KDYP
rQXj1R4/BDtfu8JcWZ45CX9TuSB5f+mJOezSXsXuDvreleteELhTS+F/IgTisRiih7vkJKUrAaIj
C5ESdluUZJV+Kkpu7oslHTFw58jVl/DtE01MTNXHPZ/JUZV7joWxFB66dTknQm6INIddPxuJzbkI
B6CnPrCjFgARVVKb9mUrzD/kkbCTr233GxYwx4YQpU+d2I/aBqDikagDnMaiSOBfOZS6G00/LRpD
OxaH33nEJQogkCG9zMx+RjfEfdcRddCrbhpKhCpxgUlPpsLkQ5op0B6w4noJ07SakfBZgkWTugSa
wTY+vfnP5yUPdnNNuTrm6SNoMING0vC2uT/x9ShxOUFJNpOLcQ2mQb9gzr9XMRC+kbtR5QlsMBoC
pbJqSeq8ozvXkV6fGNJqctBQB67nZ64bruzi7o8c1dkdma4b97YtPyzo+c3LZzlowEgCnuAm0n/V
9e/pm5ptJ6x6yl/86AA5J7srf4IUO6zo/dy5PZscfLFKEK/w52w2W4V81G8hpWBWtFgkD9r3Ad81
DSOxfLJ3Gj3sZE992pzBpFw/+Z3Bq5WNmOQnK83GbIy7qXnIYLq1FHIXH3N6uzaSMKCLnxSH5mPU
wtWtakgfz3S4uZAYVb1hW3kE/ecRuW7x6WYzAAkiKp+WH6DO5XIcGG58yxdvCtSB9pKayyQ9w8D0
qGJmy6OwBC+eUMqxU868YUTAx3Ja0LJWBub1kQ5gBB3XWNfWlTSNW4MBvX6Csccl73q7JZ3YdsJF
5fLIEVJeFL8wWM7BssYkafIttQYj60XF9b8Z0Xm4kMquSJQn4LYjawcsud+Nfrus02y1BY+DxR/n
dHWnFjAHS24+PSelphmm8KgMCfWW7M7M3Y02Xz7HeqXzCV6pP076xZTBew/ULgs5uZrsEgVbH9W9
cjjzgJqymb9D/g5Qkg6oSlOMm7c02jKt7TOO5ETgjFkcQwecdWvIjHBWPy9jp2xIS9V6FkOOIYOx
ZBt3HEaFEDLeyyshCNUxfFk31dhPObMJql71eYXVTgv8o/uy7B/WzM/yNSqzlqCrK+l4d+FoVDxx
HYLmTzkpGTtnDLx3GRRDL0r9SZGNy3YRUWSSzWMGaNOP+U5lw+lggmHVlyqIi7p1y8PNmkw1jsXp
cAUZkKkTg8RYTxrWY1dNq3boDQsuTGs7j+AQN/ED/REE3IVbGR8zNw0Im0xpoEDPI5gxsjk/N1cU
sjTOexXLMs+8MNi6qvUNxJIiq8l/RSzj+x78FL+O1FIf+GcwM8X+XblyaM4lndxHCACUKB+u3HW0
TRAPrFLOh06ZFv3ugeTc0B9DZJLlI8b5B1k3clE6+I8S03ktTYuu2LPFZ2KawygaF8sLMCLr4ASt
waR//UAZVWgFOX7J0unsIpq6qZTUIpIWruXLasAyTK9PJPHcfQbIxKmP102aRzEYNO3JUK+xCOey
owANa4J8jugsCP2rjIldDpzvMXJXXl8ORUICzFRohOGxxe9OOXsEO9hzyhUO4sWlweHeZVFTpL/U
9jK4itgQZC3i698dgS8fY/IDO1aSag1V52rz+oXFj8f4vDHw8mPfxuPqGX0KzqgnABTFCSb91d/Q
Pa92jGaL73Ent83/6oTvO9SDxx1En0qGQMOiTa3ykiGcMqcJf4PPT0VsUbXSSNXamQuhT+hxmAEY
/Wj3shf4rMoyZX7l6zpLP/04J3PMYo50/+T1q6WqDAJlKuATDnyUhubY8M7p4+iyiCbfzDmjhmNt
bC53gxL4A8tur4k4E9bhU0HBNh9MrHgNrgOESU0cKhbSHnVieO8VVKK+BvM5UYjmmEehmeXGjE/Y
3aDtO6xmvSxfIEfq3Z79hhUN8jeF8fkElCvbTO56kE2ypSCONCBitXuk9LHl5MLaSA4rFSdtspzZ
3JrO9KehPgUtt0vKgcMWp6Cez3oxYQTEkTf0A239vwD6V0G49wCuh0Fn5dek+uPutLUZw6kIzQPC
ANHfLieig2e+GmloNlnkYyq0i1zKqeqF6RN7bZAGTf5EXNYC6AK+QWDCj0mLDtBkeO2bDhsQPlPl
LmI0h01ym2iStNSJs7Y5FQoq3PFgT5BR7wNW16aUOd0cyFaQvRYkyoX9j7uRh4YVlvr4PBDQQn/V
+V+cSAw+R/do27fCVhWudJSQAiJvJ8dqOIZyoD9MFdk80hx7aLhlwhGirBQSG2qSnXMiWAiHDJ1W
G4PhV9UfsMIOFcT+gI8jcnljlUvxDPg+YcRGR4bOieGotRlo9vxJSo/yzWQu93D3Jjy9qQlILreq
VRpmCADM6hEkj1amtHp5cDYSTXMDokiY9J8ZYZmYBoCjRB9B/kskxKgmPuxxcC1v3hj8GtXYMecu
+o0Aw+GOQNcfiDwifqO5nnW4+EG6PEXSAqtansAX2cPgD283aqdU5sSWiOdr1PgtU8U4TunOgtNA
ZsLodEdoxhmGkLKpPpuZzHzndxUSlVdpInAIPOEZmRSMToXer48CdBcYK2mFxRT0ZxfuGLsUhGGk
k4/81fAB32HIpw7G9vH/wsfaegKcFjen+qbYJF0VUxwyfiEXkRWZ4II3EO7ExaLOy6gDqQeFLntY
hK6+ZbwHLzkwLHUR2blTYXO2k4UpQV0eIakk8aJ3HG/qeqF7/0nhg4jyzOYvlWRi3piSJdFUj/eO
0Te5p120GplosNlsgAL5q+wqExLjP3+RQA3fy5Sq0b7oOhNTijzb8c/y53f6q10T+vOZO2fPiSsu
9S26Oe7gswd8MEh9FCFpI7uQvB+LcTSRYEHWkSLXEIK9ASB+Cp0AnMERoMDqXIYFA2WOUw46kD0H
CLPibgqVntS60q2DRd0pICf/lue9Q4h/hqS2MEr5KrChKd5VB3ZIu6Cg/uJV73pon3+kHbxeM2hu
JsoUgAxU29s8bLXyFQfVXO7Ok97wDyYvsbfzWq3Laje/ru1R6P8Ub/j00fk/FTh/6qLDUd//iOw7
wxbTj8J3jaZN82z2eg22FxzTJZW3HrTzeanJoN4HgZb+nKYLD20e9oKbvmdPSURm7vpagHyNYYRW
bEEiZxrIXEjLYmdLCKamlM+Nlf681cQ6crN1b1QHVF/1BEQ1dDZFV5WsXuIB+KMGbqOA5kcpvu1/
fRp7GtncO5VpnaA6OpIYZ8tDEkSpQOjtZUVLztdTezLqJp+ryoRt4Fr2nmwiMjRZ7UDt6YthAXRW
uMBZEh95DZQSXP8WkCtPZN9Ye5iRF1GtXhuruIUL5CETI7UQ7he+kLOZXvqdepeip12f9OHkaOdZ
9ONDvFzHwODub01ueg18OQ3HFLIfbtzApj3yLrT9uCWlSdTLyis+Z01oxLTpbVvxerfsak95WVOU
Uz75m/S2+dYBFNmsV9lwc+qWtIDRPfcmP9OB9nkH3/p82YdtDrMnbhzNV9MC/UXnW5IqIL9dKGB4
wyVrKgx7pbscr9If81rpv9AoI+DUu6Mzv+nR9wj7yCHbqe09O9ZW7lnM3Xx38J+UqXjCyYEOIQkk
HqsvhSjaCiVGptGGUxUPkS4OBL4sIYNjavOp1iuGDu7sY48D9xVZVuRKh9d1dgpG9UFFw4TuqwEe
Cd4mMW7DjoBA59RtxADZx0maFzPKWfV4HCxSR1DlXIpmP1Vlzkf5TrFSyCGuDGhLjGsoWJzBGiVz
pcgjviIqyt8wEaJKbIwGa0w7mqxUMaZ+qurjdNO2el+VfAbXFg306Q7jlcrIwhGLIsnI4lFQ31Vo
boPeBS3ctKvbXNb1X9QNx93j6sWqtrcZzRQuJKkVgVeltXxn8lrreoqPdYRoFRiH0MvBd+V4GWL9
9crUB7Oy4DmupyfLWGsRj0S/vt5GmIml6QMstJD93XT/Xc3Z/F7bwaqfZ2eD246c9quq/Dj2rDg4
6sl0B1lPbBCq447EpBKXudMgHzQEHENzNTAymGaxzCxhGxY9JfqIgmPDsFirGBsWz+oPGBg9+ODh
kvtJoMRg5GmHs4SyPeCPsP2HVQ/oU3260fYsWmHE3VpVl64eSUx4pCmd98byEOepGBH52VZx/rJR
O5xp5KrnO2h+1UqWiWz+Vip3sqlzi3nRz4nSZQFAVXKUOkvLCBOYkqY6ha8je90LE2plxFg5ob0N
QvMYrJd8guGS/1LnJDGqu69ZkvijWlFYzBEWjJRqvWwyabyukmlMiCXqMhQZDd6LNGP/M7lY7Pmt
+0Y0slcH1ET29aGHsOHwcqTNZo62z7GallT7h3y6xJm7aBkrgKgq1AZk4RzI5BjoSfoBiCeXdYiP
Z7ejhj9D8UW7JfsksKbPnh5g1F7Z+ePpjJnjB/DxVNmaNyyTUGjR9TqBUIX4WTdgMtKta8hfDlRR
HMpnmkPKeIlf92KOBGmQyu7Kw2PFVKfj0u5scq6/V7ISzTH3tAzccHjP2WhAWb4HFor9/gGqAtdp
+VCUgypLWvL1e/RRmVOxDBFrzO42+hO1jqGha5wh6/bhRRkC5271joXvKKli7WVtl9FTOc3lDWGH
skOyVN6D5enl97hpscWXIlJ4XXBvyCFvPJApcTBPfHI0RNjgN6mg3RvtYQ1VVioT4GdvmzV3l7dP
sJZj4ha3IBCfJJvSYaQdORyvOuEl1OnBIK1w7vxwJseTduPm8FdhuI8sbu0W4ZdFs2v2j6/5YdIj
OAnt9HO8PCJf8b4n0jKe1a2iiJmY1VqbK8M5q855Gvw3FE/64LmMF7lUCBXgEw2xkNd0lqExat1D
A3QcAE5kzcRVmIUH0mwMG2IfWjOzp0dag+QmIsZY+KZX6pLjDZluk8L7Mu0heq5ePDresLnuMZbZ
q2Y/ZQTEiMyN53DKbPlt7XKQT7GHpRCwUykgxIRagllbTTt8aVjbPPsS9cxscCUCcQvXlwfVPA2N
M88mBTB2Uu6WfXbRWxgtbqXoD4ac/uBSkWa9pCECSFxBGYWczx5qlX99EKgAjfkrzGg+nJWSKeyZ
jgSQS8oRU+8rb2EritpumlKImveS1zgANNXOh7UOxTTlKIAFnyAl6OYFP6wEYvknkelGfOd9KWRL
bF19snQhq4IzDDc84JGiY+Fe7gWky+5tLINrVMDMLS9MbVE4NodCpcy2MYOMAgHs7PAt95ITs1Ys
IKj6sNRPTZ0yExaDSpaYvYBbnhH6H0Be28VTunBEPk27cBAY883uFx9LH7b+sVXzUqLRSH8X8bgZ
bSU4uCvZUIeoHC5zdO94F5JAgr7Y1I5NZ5VVR3pWGaA8yl6orkjFOJVGM3B0X/B58GQzMGvHNHLw
Ht2Ii0Hgs8leD1UtTBlCamwrzZjktOAwUXlEUFaIr86loMtY0hLel8PqH38eZm8bu9Qszlh0/5c5
9jm6Qz5sOLGdjsXNrxzXCLo7/dmPqR7KYCIq7ghvlXohJbr9flB5T5he3g+Fjv/c0aEhifiRPPni
9x/uKiS7uslcz2o4oQylbNWCSIHJXIRob1nE4aqk9dGCgrVzqv9cNqnRrRnenl5ozeVDyvTzC2WV
r1xq0zPi1FLDuzUTEF7qz5yZe2cy7pzsb85SoyuvnvWCZspDvbZR0aq/nq6+sCuyFh9kb3eHgBet
lFUXvkTuX+bo/HRpuSwkmHtZwTYoRfk5eQWCcStFFCav5YyOVj4c/ySUi74K7E3S2s7JvCTOZDFS
gSlY3xm1ItwZMrAajlgBTVhkbWZ8rOWc+W4GaflrBcXRofw5GZxfMVXVYXIxYo+V3X7ho51m/E5+
7V/39V7IThmdT845VXvjM++bXHp/xg31dr7uJdgunlGWPfU6Qj3tkGDD5vvqXWytzj93GrptzDX1
00T1oSRl5aQiII25MF5i+8qhlSAme7tdC/dAPQ5lsoSFCrJFst0n0W4/e99KbSTqnBIXJvA1aY5l
SQXvzid6re2UrOvx9HRbSIvjInM13Yrj1FPHpFU3elYFyhOb6xkSMDG5vRPXOuyNqAlwS8Hwki0e
Rlrfihfl8vGP5YNgow9gf7fA4ThU/kzM3Re3E81IkZrRzHjJ0vX0BTtlRq1j1rg6NwkhbmmadAW2
1KiVaa3FJN9cmljxquEsoeSm9ji4ybQ5gOri3MzgmkdCMiTDLKjbf42RWcRFJZwCSooJkQ/Jh4Nr
Vikigjy32zY7ULHkA6wLEGXAqd+/i1deKltd5Kx8BMLFtxkhW/7TfO/Rp5ebpfY3py06umc31hcS
e8PnDMRgdvvXyp407nggvbMysvW8nqTLiYo0tx5+OHOZ3TQomo1EBnm/gs/WySDiTMB/IjIY9lJu
01t715C6FDBrJG4787RG6tb0HcV1LEwqBHub4vuuGurbdiqUEbuCpX1fsYt6V1aZIlnO9paQUrDc
+AzZoapqAsy514F9yzIYiViedkKFrGpD3JumI97gZx7AIbGH7REymxUW7S0KZVNzxiJortniD4yM
8fUm4pWBcB1BbdYyTGECqeat+IccZZ0Gr5lFOpWHngY3AR48UBYmIUwqAvKlYn1OjmkmdlBb/ic5
t2XvJVQuUG8M8dz/mfNZA3pVM0eG/bg4XgKl3j8WXINT9ZVC2OiJwPYgFlUA9TF1C7l5xYqj2JDg
h4/OAEgkrfn/NQn+uc4UGz+I7YPYJmrRKsQJlZmfTR818FTiYkTZ2WC0adcWdBb1ilwkukCFlAcs
VZWzktcDfo3UAzSPgLUX8FUowZDKHeyn/zkR/f5FcexlWaKgl7UCcDWy2FhZs5TbmwGgY/kVKZTu
n2IHFyJJ7jq1f8A/MS3FlFhN63UFh16PFqg6pDh2CcyNbJUmOCp6JzAJVFAO+FaEG1YOG91HVsGq
7dhUG84DvJFJD88O6V0/eDqIeibaAYcjM8IZq72AIngW7aXLHoGiyN1/RMJXC0aeL0KF7ceqvXgt
c5YzYYW+6hcf8KHRmXEfV8uMLS0fllhAHUIth3Lh+pY2i+uG3r06qi5epYz5h2YR3OzaGUKnTvWY
2Hp03N9ABxmi8w+0G6GOMsrz6SEJcR6h/M9p73WhhaAkJMlUdFNEiufliwIR99SScmxqhEtzhlHW
4j/QRFHfpQ3lymkQfkVI6gEFBk0FcBDMkDwTzoMWA4NdvZWazz0RunJN1GH7cj01JYW12neJUs5m
ZlkndSBMkJWqjQaUlKMa6syvKpnCQHvAFR47F2I7UVdN9VKSJDjqKv4uPiA8zmK5aCMcegR3YmUb
HKXbAGoysw4PfpcgTLnGwzzt4n71FsFQieVUPqm30uaAjameCvJybSrQZAbcCQBEScq49VMiJEfm
HaXCbDUliG6aNRw2Jg0JVTmv0sVA5SmkcKSgY2Lhibl1eq58V5befD1L0OBoakO5AzVq/6/6Kakp
tB+33O8eYtF97TW9OM/tlfwnmGYyWk+1mVDdTSXTf0bEFjucBjVa1bQsKpycbqfNJp6V4u9S+b/X
JPmLPNvz+Y2buHB3BSYa9e8KobNR/hp8ra4TSHpw8SR1jtuEmnZ0RFCnSVpHI4cT2IpzvSf3kvqI
xx6Uqo9Xx5+lUjf+58E6W8Jc4QAYFGMckVMr+H6Z1nlhtNhuoNPHtyzpb/o7yUXv7+X4qbKOmuEK
4v6xeOTS/+f2qUPJSX9dTOW/BHKqRRDShd/NLnNlTnA2tgwVM3l5VJoLbOMnPl1M+0Z8qcIh9tnn
R7UQRgzDP0sX54mO0fsX0aZhOBeciAtjvPq8N8ZtXYJlS9q+CX0B6uxO0bceg9T4Fc0WKNAoc6+4
GJ90d+WJcWuALHm+TAtSNz2xivTg/wOn8FBeFDPv814onthiot1AH2+CqunJPNMHdL7lYByvHeVX
vrX1szUXoLDuhUCL1sLbP4UdQh/+PVVVLIMAHdl/QT5uwewN9LT+evK+3CUOgOLcTTovaMS8XQ7Q
LlXTZjR5mFgibLobkn+mz6lvBCCYqMtnbEv6FLf9pkcE9iZKBDdniM3uvC/bmEugrvn5HNlxoBmH
0kJ01LTz5T0EuEDbfav6UTuzdeH+aBEy3InQXAe+67+A/TtIFVUHCikbVD9RvTFmibODLHGNjBL5
33fkwTgTn7RlA4RN6Jdc1PbCOI6QEpvrGXrsVjyBjL2WkRltkqLZ7oYMFMad5xOqo7jX9Y3hsHza
gW4BjXcFK2pL6lY6jV1n8Xwipru9BEkfKNAN0FI01PvNPxII4EqhrCEfPPg34jSLf7JqD1pkSpXO
oCb8/IbFpP7B/jJq+p/MI9yKmjEO9OCMV1B5HdIgi4hmt+rV6CkoUXRsvpny4zKfgJxFivhQj/gU
ybo74Kwkj1PePrSReOdvEpXZkuhbi6f4L0V2P+Vg1vjLUErFjsA8Tzt7r9ieCclhGw1hV2pbobBp
g3MoiWTqFNv19MN7BoWbqVWVnA8xj7KoUs9XFPYUkxd53DoeC4FcjCA0TnHLSa/ZEXxuxnupVKcV
tphFNgm5Rl29Ots6D6uaMrmfj5nFAiBFxL/t7E48G0j7f5HWyz+boX1cLbdybz6hg5NEssHQI6Nx
wPSHa+8taiqxQA3DsgfkIUMFq+uqSIcb8yA3WvMIyxHslpampKnuNWHSnNrm4QdylAn9J9chdZPU
ei7IuheN3PBqXLa0wks98rTktxitcl3Pk0kZmVPnQN33LsJnFDnlizIceGp2k0KXSmcz7CLHviLA
SM7d94BNCso/Hr++f2idKD/2SsvVV7ebpaFHKIrPj2M5NBXV3hcf3RO+EdCnddBr9iTAlPBJo/1n
/Ww7gQS7KCaokKoJ4oR6g0LrKZDeSQTaszGsNfzedd2JVcT8nYTbIoQEwHfG+t0/0p6+7/wZ4MjK
RrHWwHcxJVi3Rr2kMHOhz3LKjaor0ZibupvkrVOKIQDc9IL7he5ug1Kj5e2ESoG096eW3DCMViGB
4tIbEGeWp0MfzW4YUPmuZ+JkJC0cXltq30BTeAd9xYv+SH76A6ZBJ4YGadAuIa/gR4uCJZrQOfXC
eoDnMWFpm0+tLXffHzqY4QmF9I7+5YWnB+c2404fCPUB8vwtW9fDxY5Ob8+b1lbL8MEDyrXs5qq5
/C6YI/pfxrqvN4vPpxPp5TGT3a7ffE7blKTqxh8UbRn/KHeNpKAprx9EPzx0o0DXKfV9tg+UPe1Y
ghJsIJWyvgGut3a6aWulBBhZKszLyaZHbRETp/wXyJ6gZLUza6e0U4sKB5CKtdWiWZYzuQDb3jhO
KV2idHGl9gcF7sgOJWIMkUTB1Pd2N9sP9oXc+5edykeezK72iXD3XvtkraWzWzCwj60uOICiNkmY
I4OHB4WK4+zhbGR6coEak8Ez2nDPfQFJs/lzu+dK4RtBw5RSubI5rzfu9mO2uvoHdDPKICQQdLvP
rBSL8FZGpdYKR1QYIuL/8+C7s2eIbKR6RpGPQItE2ymHfuXQrFKKhPg5K8S24HfkiJKvD/94YiDX
Q56oGSnOmrn3wGIATJE1Go2Kn9WiE7wAKctMqXfPTiUwdzvqbR1XzfwGSFDGXgB3Mz+wTFcC/MuO
1Yr1bAb2bOzGGOTSKBS2/rRvmwWl0P2zbgRSpHoSPfULBE/1VS3mcT4llzUKS1uj7v8+9At+A8qz
kWdxtdLiHX6WJ4S3QZxE0vMjQ1eOHuAfchDcLSv7w5qaY6XrdEXOE4r3BBs7AqUCBecOU+2rotRw
Nhd7I2ZZ3IoAFI51LNAyIrMgEIWdpN8gw2ME5PhmtJZHJLIm9HCsRtjGOjGTyw5+to4ygvM4JLJC
PtDsOppsCMbMN5gqzZxXHZyFTr92qgJsthIer8mlFLxNOnT17NebWnJfu/t7+rAntbpUC0sCIwx0
bk6K8Ol1iry+6HFJB6ctsPz3ZsUHo2/r4vokgOjimEv4ec6w/wNAcpCNdQ6zsx/6mWhGC/6xGSes
U+sXja5oSXafTSQ8rMtTYH9TQQVvTC/BVFa12WGeaLOgsVwsGYp/v9QnYqbTA4z02pokRL/wFoOW
VkkQ1Su1VX5SCVUgEx/uyMKEufYoi5HM+Ek4aapKWqYxR71+HaD8vT/ZiknOSB95Xyt/BUWroP8S
frLGfsU94I4TanMkCOE/R4h65rVqWefN6sMaElfYFY9GU/kE9Ak5sFL0S+BB18cbkHEOW+c/8hwN
wTuzPGvVN8lGWLkz+r9Cg9W8TLqF8Q+FbhdJkAw2HzjlviJdViHxhe4z6HT+FoFWYgJPWQdvwKTU
6PEqw8DmFiGj20UOhU8DGx7vIqbOh6Fd2TZqjySHLLSc8LQMCdETMjDlTYBRcHrm+oWC4Vo+kMS1
4sfTT7NkL+c9ZPLvAj418z5V4ObL9Lw86wcFM7AOzAUFHbwob3P8IpVYqjxz6N8CB6gTJXcpWuIj
wbWbkA9J4CeKFLYTfzsdMgY1DMkDH0vImLGmUCgt/Z6IVAV7m4HaKrIm41egDlsJ6fLO1XkOZBjG
X9oW5Z3DOPBky1jVvZa4Qht3NJ1SXj6zexRoJT9cQcpyBd8xWJwcN95AfQmlV/rZq9SWruX/S28m
SbI1EHCBUspeL8h1jKfbbrx7bzNWd5UcVTeBNvDt5ZoHqt94UgTjO742+RC+x41x9nRdlwYsmPA0
P7NYldiPIw+g2t0ki3vzCi8FB3E4YitMmA61zYJETa4hySOjCBU4AWxNX8t034QKy+yybmkQ90GP
dNzdhT+Y738Aw/xNVRm9BhKpjc75B097VbFROlzPF8xKZIbnNCSqyKjU5phRyKW8ZDk0hO2U2BXr
4gBr9kOay1NXy5QyWqJl4mCmLVJ6NRerfIAjNE/ezRO492m4EWZN/xP5JKLycV2uIzc0341cfWs2
VZe4JTrzZx7ys8DcSasAIcj3b9T5qn22TluZBw+jk8R0KddVL+8kkBS1UERLx0L+0m85T7goiX3q
jt8ienWfDsvJC21t3+YC2LSw07lM7TC8npEgJim9EOJ+Q8+3+R9QsBYeaE9b+N8YTUb72KX/vQCr
D7X/VARp+2IeABNvemGIt1XZ8RAtK9Boc3V2qKxxJR3U/CQ4hzwXvQH2Q/JeNu8jppDFJlVrqhV2
pFGKdw0Ar4AudOKpdILWWvMDDH1iXCMeWdcNLSfKP8I9FTaCa2xE2TBgg7Z2LL+NuFbZ6kXCTcNM
14y9ZoFQr+hpZjBCZf3e9otd8V3QRz236YF7afdeadEfUP80cnaOTybRwt3zzU+10ZQqI7Y6g+WL
o9yCF4JTnQi7bYWxWlFevp5OW45TTY5gL4uGvqIx4TRNoFc+94l0dxljfOB8y3xzShCXTIVzO1QN
RdnoY9ay7qlrzUF+zd92xDR+xiLLndpRr7quJk6Zzz6uDIEJ+umtwbiplXvFQVjb6RQtaevPVl/u
U3VtTs///Wh7YUbCTD9HcyCaHtLHGw6Ku5T4ncPKuVuW+sJhnEFQzRF1qYODAhbBdhu1hRbzg315
wRXLT6n2aICqWvoR2zRAAJpoVs1gJFGdJSmW9HzCQ5x08XXaVj8JFGJFbvKyjAaRIYJ5KYALqufU
KFwer7g6HVIeCrX4aolWsjyjyXx3D9KGY2JhqjWWHmQd69P0WkdkwKC6YnBNQjPOb+FuZukKQXyh
XhTiU0jacI+rymA5lW3egMsT07jHddBnSueKdK5UVdKVzXPlJmwoGxzKOfWUyc4pVIGxeKRjLuKP
Uo4KLxtojpfJacaF8f1NDmESjbWvRNPmnVoKGuq35iyN/3Zd1UCIlU6KGvezMPIwpyii1F2/U1l0
7mfoDoTYNYz7HqyVO7VC68qKgvAlyv2bizo8ggh7jf8EPwPxKqTgWCLRhWteA6q4jonXL+hQszf0
nDdRgti/udC1y+Z2E50K9WrAbq1YtFVg1FuTKePk88NzXUf2Z1nWxU7HYbx09syZDiJ2RAyKEv3b
mI3Zx5iMQE3JKDSnc39rwvS7VkN9BrqAwNTit+TI00Kf/C3T9r2LL2xKEqZ6dBiS6n8R+3YmsGCu
JVxiVHc5MkDdC51yjoApkKva1FZ4fqNRk91eEOWrEPh2LG4DhRtaDVx9MIjV6OLEkDl7DCuOpL20
lae+ge5/Qw4JbR8ognT5t4qYY56aXTXsu3llhnwEIV/rabnhrTOiLtVg0kPb42vvPcwlgPELNU+G
NkLNXJAsbts+E7crEOgs9CZIGZWBgHVb3ptX+FPuCgVKd/RcX9n8dZMfvlR0nsOyobO1HzImcWvJ
oIfvYVGwTSnCcmcmQ9UG3OV2IfrJg4NpJTgqoxkoHzUG/CPtUTAW5/EiejF5pO9Dx+6uHMtHsc1E
i8rKYyGfgG2bb67qUbm4W6Rf3bkyczf9zM1zV4EGFtZtMCSMccRZNVP0q6W94pw8p1697f1Dn+Tn
MAnDkNPV83rxyI1jrWi2kvZYXl83y0tIb4SFySoTBs4IG+aV13cORn7cG2QeKopcu1DMVlWtsS4J
H/V5KStrdD8ZHwyqlDCyEpfAqPpCK+uTukIbd+3zTdvH4udUsOIDjuqZQp8doQFdSoaV/IiR0df9
aNeI18Ma4tF3sP33KgTvEuBoz8PgojZb7CjISUp2QCPcaQMs5EJWZTHbaW0YDzfzKT8mi4vD0E45
ydan3GotdEGPhQOq2pJVpYMnEdMgXWWmWejE2i4r/j1YeswMCywdqQflxZtA8OEalLJ/u7s4i4e9
iTyuzDGL3Xzs/FjZju3YEt/+teAph750pji3HgmYdTl5JvHFA76zTm03lTHE4fWZrtq/lYJzFP95
ZknJVdkZWbazN9Sm20VQvl53kN9oiPayLh13ACRr0vma9K5sWrDSz+3uHF78wpjf3QvL2aXHTtAz
J5Dy9ZecHeIM6x61iauXwwPphGl4G3THlpMJMIdyXPLy1kxkqXOMd7EEy7kCj6nViG8kXBFxEstl
YI7Bqxp4lF0BVlzQMesO1ZBcbb3NkcedMFJpCcmCC1AcIaIBfkk+EKtj6esPrTdi7y5PmoHAzkyO
LZxIbIVGONk6PSTyb9q7zPo0tdFGt/F1q+as7FUF7peQkOIOtN/IQCZ99/YnlgE62WfFH91BAZrv
IE2ouqDrQYmNRuflXCU7huKrBCUo1bKiEYdHTmKlny1/MQr+IJRCI58A+q5sroYJQ0//EaWch6BP
0EwijHIOBE0GuhR7XwwqM9z7n723TZ//gYXy0uhv0YAbN0iUYoExvY4627xqixTRlzetvg3RjT3N
iiYHPTwvBRr6OeZ6Tjt0jWh/kiDXYC8UXg7E3jNFEEKYQGnPWUSMiHr42KH7kTBFTwDakUptBTAY
/l2WX2GjHyQ69b8QMstoInivA5kBaCNK/YDyWCUjeZ6jfA5XzFKqX0tgOpJL9i1QNOv1MsRD7igg
yGcimiJnpekmasPenuAxy89umGc9v5JVHapOmdgODzDVuAf4oFQLN536734cwjF/6uk/r3hzIapn
7TN17lxV31qN7lS7XlGBV2zPQ2oVToQWe+HruSAKhEsl8ShEOhUHYcHAN+KRxlQOFvAtf7/mYJwU
R42jbQFQbowUwEI7zkuTvCNxLie6WN8eFKT9VjJuEAPxWcY9QIFjpGH635Cs1up9KZsJEWE4JwAA
qP4JsT/pXrsBXjOVuXtjHwXTkGxXB1HcQ3qGTbKxm9zalS9iBZr6/lDHtG0++k2v4RQZ5sCD7rKu
T0RyTuxZDaU+T0NVVFNe/jyJg/K1nRxMklCEQoVbsLxBVa7t8gh0Ua7AP0Z/xLpuDY5VfnQp13L/
83KoUJp5V7dLTBRKrBm4oefmgzMoxWPwzDXmZnn900W7UOJKc0DyiO81GWXHKBiYvqoa0nG2Ok4R
/kRuB7UnuM/nioCjiCcGiEwF5yBokk9/bRsDNOsdQD6nk22L0D+9Vg1PKwxgEZ9EUds5zgVV5np4
9cV12+72AviZxLQovh6NEPd8/MkFGQb4iaRQgl04CeFRAssO8CZfW0PsrRD7MdwMcI//RRadwjjW
k2N25mr+SaNLLi8/aANHffjCw3bj6GaKCRUY0ycIFpU7o5tgsNbQwXvEQCkYXMvW7YeWyWHVzxqJ
RaOy/KyhHjidP69OMUF/BmcDld+dsTILixi9IAQXVhBbfoQuBC7mcAPvLxXOBmMiJr16CLfg6RWN
dgQ12DZ3wYlYyum9zcgUTH002UyQdzOyLWSDyR5J9DmcsGZapDYcr29vJ48rxYS+4HJhLeufLLRs
21nn9SOwQ5bJLl1s7K+goCa5C8hpjQr/KfdHadu1jQl//dzJ43PP5jwNWubIpJJb5oYQA12pmrcZ
GHoFFY5lG3le8fV8fhifRujEk4ZT7Yv5taeEc0bAxisNSz1wLiN/E8dBiPwXpdxIlQrv6MZxaDFE
Z92RhoyrJcflM6fnayiqHbEKWC/QX/q4Y98sBeOCSF07hBiqLiuRiJiyRIcrfJRn0DbGLtzlM1du
p7RNsbYiCFgAtemjuBEJ9eUj84KIo0d71NFeVBO4tNTi7JEd35zHjoIze8AKthCxfF1LM37OT5ef
yCj9bKeYu3GeE89+ktoSnvUbC62jlg13xHidue3Gru4cjGUCySp++XODrwcHuxGj+eIT4Co391Xn
fUiFjTXXUX4aiOPT0x6n832UOpnng+0yzDsca1pZHFNMaIES3KMHzbi29gSgWyrL6QPIlk18y7x5
+JYA9QNjL8N2Xcev6nskcF/GWn0P/n53wNqhK1R3Rhz4JqoBMhPuf8/eXx1HqaTWexuWrbj0SjRR
29pI6ufOBH5YBmkyPoOoXvq9DEAbk0uCC/Db+XBjzIPvwXME7CNBHPaHTQzWvNGXs5Hm1O+fdAVn
ES2WROY02ENkWxVh/dslH45zX+nrlaTXEgIdym2ZeBx6Q5QBdpRGHI78lQGC3z8i63v+675CTZ+I
AHyjqYqBBB23VQGhEBYmD/FlHTFpFR6UbSQ1LdY3SeO3sDsMrMhgt8JOPgeqdiKpOnsY9m24dQRy
R8P1AiCvHVkkMG/xCyOvg+gXZvVLowrdL0XBF/gbTrOLIUnhDoz7NLwPYeVs9as9N77CzfSUlJhW
JiZDxe5YFuQDiNNeBXBuwHs9D2sTXduOZdrAtVa7Zb10wR9BrI4tCycdek86YbH9++6QlYlDYKSK
/5GGgTIzMg0F0VOcFhgnbAvHUbo8Qoa8uWZlyObvYLt8NVI6qxI9qu48DJOrMUIlxDMxEiqLyo2V
v4siMjBo0pho762SQWDLLIqrSr+ro2vHWxJxEguvzVe2vhkdDF7cab9kN4+lHhIjnrwduUKXF6iK
DNmkqILhTb3zuy+hSN24I+UGaHq4AizmczImXFFvVefB487Gib2EI7LQsaEKwaD2StQA+QDK9znf
S9e4hRbFDZsjEGRHuVVuH3Qd9+3vbXEaKYm/HrP3B9Mkvr9X1GG/gd7ITPm1fn/NxlpwnmUs+K1s
YTZT0Pb2fa59uHd6gOGxx62OGopY6Cv3bOrFJ27kDn5Y3CTjrMs/wbW+PgLCLseQ/r1L+SNcOqKi
pDQzzeMEG5YuKanRDM/X0lZIe40o4dD2g+iDNUNbflywk6JFMZLDr4dnnAxD6xsDCKaRNpvgFYOw
uNcwDfGcHQjtcHv3EyzmBtwnKUAHxWcET/d4FN/Mu50/DWRYSHxh+zUT6yuAkEDW0QMyGb4jdWzT
EAB5ESiCyoDcEz4SkNI861JVLIFk694Q/uR1Vr9fj+Lyj+6LsP3BojIQKOb5rjw9CwLvLdwulC0n
jaKzFC/FTkgglfyB9nKvL95VVtSrdpSiqL+SsX3CZbDdkCIuf4mTRDT3B+SUWyG6KfQXnkFn14h/
yykc4Nh9ybOzsFIO2QEQm12P0NKgKCrezCTjyl36LJxyFnY4THIlCbuWYpK2i6L4H0ugVMbiOXvD
XYiW0kZuO9HfTArcug4VAesbtuj2gQBRdBimvdBqFzlyXqHrFSb8Tevhe6KVj0GxYEQUpAKhjoSY
tqTh/Fany+BfrX/FbWutIBukWXY2HAbp6GEh/r69IHG/S9VCLzrwveGAKonX2lOJZxwjsdNiLyC1
GkNmD+lFLCNQW8VzOL7qSym9c2B8XP1UV4xORT/+Yw/yImfDpO3EDys2aZZsqyjoCzCr/m/ToNOM
aeokVX/O+71PmxAWGLBgoV7IGh3wpxz6SNqDQPRb2FNb0ioBSpc4miycY/1xpzImO42U30ul2Odn
2qkNXo84gS9RnOnm9n91M8+NwwghgbOhvwEMWAR7PXveydcL2mZ1LE6nFyQ7qK5Mc13i1bXTycEE
TCOlNgMwuWOfXUMijuP4OtiWMYLr2BQOGNlQYDKuXiN6uYmM8Vg3wkATM3qtHBlx4gWYsCjAejQV
Z8en/7+uiS/gzltDeNFxgYG0p37WvEJ3QNsnKtr38bkDMxbP+OrIGx0wsBh+lvwWelwSdK9wcP4q
28vgjd+1batFAlRyyaiQuaytacdofyhal6OhAvrnjzfDVWBpRJmP2qgfrhsiCDHByBc5XUJrWXym
5jXgFl+XykTriIyLj513j9SnpoHFzWPSgYY60ahyv/qHZvAorEiWcGfInYC5MQ3MSABmLJNjKFxl
ZnLT4x8AYZ3xjzq6i5Bt/hfLDlCJFxhgZoke2gfen6gvPbZEt5YA8c0ACVQWbnzoMojT4Mm2E4Ps
PQQ/7N5MrW88C4YzxmCwc628oHiYHRh6yHqO3Tzz28aIqfi0g90Ty6+10V+TdgJ1MwmCYKMLKW76
gDp8mfSo59qTmsFhyjmyABZLkt1B7CBKZoWP5wvmIA35OMORdFtl0YFb0mgmX33OiMCLcmF/qddo
LmadczNWc1Zw2ef6fY6YA/0z+ITzdeSEfhLZYIhtxgullbszYHPZSG9GwWL/kONpwA0Zvus9fXU1
fAQJcxBhyyf9AoqXrQnFiwNz/6Q27D1vVYRH3/UsRKGs4RDDPQViMa77EH9nZAjNwIJReaRVg4cm
myTQwkS5NZByeI8EtBkhwsPu7H6/tbyHxxESxGPWhzWD637nVoHJ8aonqwO2xRCbDvXFBMMx2wPV
H07KLcS7xgBdRILYYpg7SrOaKOU2XR27a1lqD7j/dhLl0npzYov4wLNhatw+hNSDI/0QGwNMsLjK
wPqmLVk5Xr0d0tLoU2y2Ozsr/r5OEgw5J/rFXnC5XqjzXSIzHhDavyvsj2TmWkVwoRlFhsbxsgg9
btL+WI2e63iFJaEE5kefKKOd+ZbAuOesfL0rF8Igsjea0bWqficZ1PAE3Gr/7i5ru1HgjoiP5GDA
Ve5r7XU15C/z+lisyec3OkJ9WR96IWs6SsT3t2g5eJT+SnpKNgpqeScexnfS8cGA6NkUR6YxByV0
LJ/YXkenAX3U9GwDb+5tNJJ1u5pKjLcLXZzGTWYSm4Q7IOyKZvkNEF937PhfsfyVyVoCJoo9WoUi
K2tJX7f5YAHMRAjGULpto0DpoJwni1PL6mCghBfkyA+3ONjCYYaW7LtitsTtCRbSmrb2FFvoEX1Q
P1nPe9CXs4BA1hbD+t7otbsje0iD795aM38Z6ObtZH08sHD6eEksbABPQGPjfUmdWwdmjjOn27oa
S3C7F8IQQcI1oNycSP9JmtyjCyL8o2ceu7meABdGlv6Nhh4NXkEmCFvTFtXCP+L6DZMVsvgatV8B
m4qk5o/BpEtQdTXRQe4SB+J66S9SSsNH13C/4WceM/6fWMDyQ1K+LgqYFaZzoKbEJpKmO8fmXxbZ
I4sO/Y2SlpDeE94tk+xu8Q93Z8xKzMQJNQmKNfyX4jdArsbR4O19akZHEOSTaNCbwEh5axMREFqJ
q/mqyWk+ALcLZWf1SK6nFZUtMD9lRQRB7sgucPjW50QQI+koWOZfhLoKspPTfV2/IqTOv/2oHd14
JfF2REPwgMNoSsThd6DZaJz7Mty3tthuE/eXbwfMNzB5bjNjrM+6ODHz+5yTBWcBCiCYjmMRv2v0
GaE2FIijGUmX7MwJoeL61HPlCMBjecCPM+8RW3MyiKA9sf9QIw+cr+5xkk9qulZJcdUgQa1FxWx3
aUfAilrrgwe0IncdDNgA6NSwsQUIBdUmiDz8XW8HLtp/OtAnGienteJZrMot57XV24/h+OsaXwxT
nF8CKk8In26nr4IaXFL6C2/+gxFD3w3gsbYdBW/ldmmVrYZoUGyT+rvOJ1biy4H8Zc+I59B2tViY
TEJV/hVcbuf2yh5Ft4jt6iRKRbZZ3024SUVW3uCnpOxmPCkWNp08ScaUfao836pVa3culbn9qTXd
85ljcbfA2ljebw9EfW+ghYNzcOKwU26+eoyUCZXZ5Q2SMXG249aA0OtZrSPaxBPo31zGBhaYdU5L
O/XtgOC+HGzqVQuXtGVhwdf+wd718Fd9/HkI1C+lJSGSlTPone/sPuh1WWJ9LpMJDZmTeK3tDgGc
Elsk29KR4eo5AttORmC5DImIO8k606hYCCKHgM29IeJijVnJcZixx4jCMuJZ2OHiANGxRag998XY
EPZ2GLC4iTsI3tJOhJ1AxrQbW/SlHN1Lbn7u2fE3rQ8Cf7pDYMu1htCdKe/SvC3EBoD2xNfvFv5Z
rcLi/HDR5fR2eXV3ww5pOok4m44rGoWXgJSD/PfV8MvOqolm2XvYMO3HqUBbf08iDSdkgejuriiL
X6r3OvpMtLdoAt5nd7zgJ/49MBZ+ketwutU/iFNZQL2ND9t/KtwMv2ZohL4TNqoZrRx6UcAHNS2C
AO25n7lHcuU728UfJ3QQwu0UIYLUfYqQA+R4CJpMoKh+NunS8Z0e3DITzB8A+A9Reo5YAR+L63yY
BWgSRiAH/n6b2iYK4wA5mT01tXX7AroQBZJov89DxQQj0pSW3fs0J4Qa2NmB+1UOYYoAQUmQmlXD
hX/3Og0Z0CVi9p0y7URYdkwKKKqJJO+rAZrzSpt7Dw3vVI42FIO0Ksj2JtV4xHtzH/ezGgI8h5iv
gVqYwHs8PnnPjgsshV8a5Bzk091+t3vTphnRPJgEyeFzEORt6mGBZJhrENK54sYdcMesFUHzmbNu
5KWfOA7sRvi2DcZdkoXwPykCV/n42JCq6H8Ps37c5rqJUqvRvlK4liuyVokIi1nMHVZWuwG0PsSj
yAiPHknWCig+lnxyv1ZC4P8dbm4TyesZro93VHA5JVl40czIUIG2eScr+k4X1gJUMNbKrbNhmXOu
9SI4IxgGQjGgL46sVqbkwLa2PbMVYRrFGLg8N07nhWacFUB2XFX7NqVRHUssInC4LuOd1IHSnQTm
cFh7ga9iK14VyNDVGJVXxSG17xzFVf7NpZWdP9MM4Ar0xDGVSOqycLaVk2mxGpmMQ8Nh+KPxRkz8
eKtWOkyxs1PZHjM4njzBtIaT0ZqyS0F5X12YtVlAhUiWUlAKeFRgg2cj4Au3OeOcxTZM6PxMkdmz
WgIBnOM0rKI/+uJhV2MIql1pDasP7/J/EXVz86g9vqhzaWQVz3ODrZNiBvAREt15TR8gxpLuGze8
+XpHig2DFCwKIcGXlKjwOFoTte8NIxYIaD5spmRQM8X9rFjnTfuX/h3Bvh0j+K/QkXzUjiuvmYVY
WoNmNiD8Ox5LAo8e4ULUMawYnGEgfaayT9tg9Qn76+vrTQWbMk16FsfX5z9lHs1cLUhFP/iBJ2H3
5+kOnpTgUm3gWdQOdG+Xwf/ad1V93HDzFPv69vzMwDPHq0mgHdWkrPBvOUu7wyCjfCe6MDaTnXAK
ybzwiDMo8xRQ4re5gzvUh00cEfViiHLOKoVf+FY0LXD1x61MXR3cJ2c8+0XMMS6O+bbnoCj17S1x
iYgfElLrBsB+fyCw+FFWDUX3ZexJN+/fASIisptfzpFpqCkHZCVz8CUQBnm3QFbbZrDXi4HSwp2x
jrc6Wym+N5ubNlCwtf0QlRbdqDxyn9zBLYCIJAGVPgy6KswxsUJ5I9EpfdB4WbIpLg7xJbi3IajJ
JKYeg7IuIKprJkynMH6ri8sym+KhdKgIpjVObkSAi938KrxWK1l7E8CeEYCBsjlGChCrDlwG+YVl
HaYmHj9C4ye9QRteJ8mby8vhS5mTLSdUzLqZVfoYqzfWWMl2FoTa0YHoJbhYFji0leP34jUiCWYi
qd98Hx4Ga8dA4+aNpSF02G31OMWHU1aQEWTRpGK59ArxtTMKTQNUVsbguyAcdwWW2xjmajUd4AZK
oUveUfOnmuVeBCvtnRHIcDkCaNuwJP6K/6QTu+DKuoS40SPtrPV++65haBN3ofCBwZTaSGsvvCSJ
4J0zwpiCankF9hhmq5OSYvLiteTaw5scVYvcsPK0OFujsCmC9jgUjAxM7lnrCCCfdHyb6Ehf7P5f
k0QxS/adXaRY+lk3VNSR8BhMeRCEDGRFQ0eW4bhfQtAV70CTEH3WVICzXsl1zDI+xNqdWwWzWIOJ
gL9wn0Zla6r9BH377RozA00JwNPzewubygH1NdhPpGeeiacfYNeYOmTQELqay2gFDSXvV/t6OIe/
6TNcjBdDsBtT+u3vxx/Qzmq6Y9sAZyIKzPfx63C6kN3WyDHe+914pOODgSRyt7GtBlhgFYCspHcP
TBUHmSTst8JAyoercyVjE2h//6uQPGJi+IxNdVnQ5gGGwprRdPMWrMcbXE9c6tqekjRnCDpjtSGO
OyXB5gX2e4I/rKcB/LM3bUrNAu0UDchttdgaZrFVBRMkm0h9EzEWgYp1pbxjEZqzhJnPlgWjEG5t
lgfIivwDd0kkBCqo+IysZ5abL7Er2IbEVl8P+og5Ro6W4bd2E5zm1lZro2laREggP0gna2mpYi9l
CeEUxQ4AmnjOHQ7EHPHrGUe2R3SRo2RfpB4gO/c3uaholxjlL/JxgeoR7YzZpS5XZ3fbb26Q59SU
oFt6v8PoneLO5R5loC3fu+cjhGLV5g9fupA0i1j4nPAuIaM6QnWcLhFUpy2lArKuHrq2Ci2yZPCp
Ua/4Yb+tQhNJWNlll7phJ1m7ibWh4p75VW/ORzYIvBe5CrrONh6AlxEp09lkRqagDcat4qIDZ9W4
s0oCWqy0NmgXWpmXiPGq64dDy0wnP1i8Q29c7nFDiZM8XOHijGaYvWyEIJfLBQiE6joK0hI9IrWs
D9VPnCW0J32Ju23mJwGUzczguvc37BR6JyrfNPGLTEbn2GcGShjaCP/GMzC07idwqmzZBwmCARCN
QIpEg7XQCwq0RiaOeSKuvtF2qJAfZkYddH4mFkdWahM93sk8nJ6k0JmjAzj91jTJ79d6jjWzEjvj
4VyGCSdL6t62v6j8CXb5vbVHSXP+ecpSaQIeNYvd8U6GxIJIb12KPLMvnrFhYgxxp16qkbJB8wPA
yTw91s0LGKQCGvaYZg8NY4wAGv2XaBkOibHWwPn8dpicKOZQanB1pxEG+mya49qzVVz0D1ZZXzBu
s++Nrt59aK8YyWFjJZz+lf6V9vQOnie8y+OR5LshSqvFQrrusDcZ6HwW0gJ25W+YhZU/2n8JSeKc
lZUlxHDF0VeaDW+65Ijj+sYNDjfFdjl3qaYSZzOwGAz59ugA3in4U8cUOWJfM9jZL2y6NajUjliO
PyCFxSCb0B//PJeKVx4tEPKhHJx8UBxkbcu31HKKh9lRYR/zGT263UQInsfuQHDUFy/iBtSuVPD8
FPvBcnmp8Gas8BmNq3/LF7RrqIQEnWKAr0izF2SBsshAEekdzrLeg21+Kldcq5BANLR8GojksL13
7kilT48NGFjpfJT8iIoP5Gsl6By/m/lZfWPmuYWOQ58y+wTXok++b078VxmyXZAT8SN2aRD+n2r0
PLx4d3X1VtxXsVLs42iAt09m930SdEAPBzGNUiEdze9bwUxiO3cduFqudemmDFFSFRJCqqmFLdIp
oJOISxBUvhvX5AGDw7ne2grR9n/33xm3gqeZca8mD2QIhHuzlSl1gP3ebDZMzvXUDmubsVGFLl0d
zscaOMPylMiwE3Q9a1zmvzb6XAgo4at33V9rfChYH8lHDMy56coO/mMthiCMy5tWHRf0U4WujKFW
9+U9PJMJMfIkXIj4uQFR1AtM0RKQTWhI53nKi8VYSB6CqzoKr/LB8aom+50At8EX/djsRLxklIFz
hpeAEkcyx0wPmLUGrmMBxYOvkTS9m04LpNVWngkHXggBG/Q4A8tS33vnmKFnDERXrOOZwkjxk1aN
gIyCux/INEPl1mwYwBT628pknLvfQXOBNkzjmVHg3VJoyOp5SkX2xhcPS6+fn6cnrTnULghuLZdH
xelzxnYvbgyMvjhAMMjQEAaRVR5MlkT+oRyuvNUDkhu9x+5iKl56xjeSh3ynPPfde1LdqxkNp1LY
GRIPEtKn/fjYnETQbMZTwz23PiBOgnm1HqijslyvASIo5iz4VvO/mBtuBr5M/YGpeoIqb7g2eEpY
eUslbrRCOsG6QT/3eJlj3QZidk6Zh6nXQ5GNKV271TqT0Dp9gAY1mUXhtuhidiY+HcRWRqz1cleD
ofMBsBNudclRxosajGmumbdqXH1m8JBYl6D4+3dRPrtoh37bseSe8r6u9a+CCFfPDJ7wkKrZGv/p
ld07uGU4h114RmFAaS67zbUYczYPyPbHa8FBHIDqGLExzf5LcksQ+RCv/teX4aybiI0ItsoaMx1O
C+1/871cVmqc4Fks5gSbQkyK2hqiPrSNfOM5eDPT51qcrkxldIX8b6autGGMfbTo2Oo4kTYTsUhT
+8i7cP45haiRnDQYJ5zrQ/t0xm6N2UBqWnFGk48k8sErVGflMeavWnSWhnkcjP4OyTqgk0ypmCiR
tY6ombA30zJJa8b1L0UVb08p9wBV1k18012p6HuiflMLaGns6WhU47QUZq3boO4yAaps9CMo968a
BDDQmmVLwRff9QKB+S+0ncFl0hVU0gADX7IEYjsVKAdkJyLnHoTVVgZy2iKKo+v9ql8xbOFtqdIq
XEajMxJGcIVdJTOx0j+VKG2Ovp04VwNLkSB6nCYfN2SRsQd762nstwjfUPQogiPGx8h5kVEGOgXt
g0gvj04k2UEeNkbmyr7TILpEtwqbWHrCDUt+FZ/mH7x20T8tJKHgdBsw/ws1FYDiW/mDwwwBAzKs
39m6JvduoKWDFsrF672dduKZs+MOi+E2jT81/YsR3NT6guAa0gsfWjWHmz5qGR1o8yumdyeWyNBs
yTWjM/KnwNS9e4MlhBdIbFOKLDAniTFB+ioULX7RDu5bIgMILIciz1WCbkgAE73kOsT1MDCVzSu7
oOaJLBKaRPPHQ7x3EKPD1of37/Nje+zIsyWSpOjAGvh9u0PVFrpKSEcuKNf7C2I1b+lqk01QuHYa
z/1gudseC34kTNiBo8oJqM2xWGhUhDvvPHl4WdpQCbYPJN1pczbZaDJm/rZqQZjvz4CdG9wnICLv
fyrRV2qsLJEQr7SiBROfMZ+Ymi9jHIB7VTGJO4Yvf65lO6Q86P9JuVqELsX7qd0IUYZw/gam8+/U
btD9KX4s3/s2U5yZwKDinUYjNyWD4PAZI3IWFp1KAWycisaBYMCaz4a/ePYqnpyWCe2XE150M5/e
LzroMQdYVp2F6qu/jfo0DSYqjTpRbfEuXvEpYPDDfRrQ+ITfRtdLPz0XMf01/bX1qj+gvxQn9lrC
xJs64FWtkN78f54vIv8f4wkiFqF/TG74vDpo3Vkwac+GCZSOBr8G5OFEOP0UQIZxTylCHi3f+4n+
Kmv/5DKZPVTDDtGEjWFd3nSXT3ugpIGms8gLu5LnLxL4OxsTTQ7DsZQ0tBED4NwKnKdh7hZ/R9ej
xcd+GPkukcMidmInxZINNhO0zXNdUPqhd9FkK9vvtH52cCeGmHKIHKp2gyVbGSmJl4LH67NbLVpq
8cMd8LZX7KgyWz9EXcExwHycFOuflIvPfxyEEDRy/nJnMqVG3+vLsDF5zbLgsIsZHWZMsOW/F0Ri
44MsgH82QOrX78vg/EfhJ7lpwKee/4lnCgfy9aGEmMOWsdgAGueQgnDFzazSPwyT3+uRS5yDtXMX
PcWze7eEAfWp8Pif8LTm9ZPKg6SRvJyidoCYVypkzEpndSXXzoCGHmbH+Zhxwv2HKAr0Va0l1gFs
Y6EG7eqwi/9J++S9djvPQazFqDXSl/j2gvvzWeRxDZoX200QDrIKMMJUthc0bhWG85/qDVrYUJim
o91fkP81I1jSm3fTDIDZGlf+XCxGVaiZ+L5DGGN/AQ9vEL5Yh7tRS+SdngOMU0NTikXFIYSZzAFz
K4cJiGRmUOFUwNUh95yJ9I2xdLUhMYTYDspZNalZvx3QKGKt8GuMxeHo+oHC0OmWzCf6pjY0lH/o
FA7rYcznKUpRCRPMlFZqykRdofCBCtzcIKzZB+el0hbdBFSx+vPOv7DAnBCoiB3PpiV6pUedYMB1
tnUJnEjdEC/HzkJEWFJKI83kpjGdEj+6weLkxZz9FaVVVuGnk7CK4Im6dYfewv8ykMPZhctpY4oZ
OsHKqJr2Hpxa9HAeSevgg83t/OVDKnd7f9OebHy1dL76a1VlEN+pTqoDbvJXnmhQj82DbFuqL9Ch
FfsWA8l3Qm3ZyCXK3z7g0D5qgYbRoEJB5RhgezBDApJzRKv7Rbe9/PXBmoB/kbiSK1dExJzkiNUJ
nu4wNQvSRpjy3Kp9Gm8eTweBnTr0fluZUPzk3DF85+rJICyFu02ol5GUM5iSDQt3g+dR+BoC/SPL
ANNdJYzwE9/aCpLSeBUqtmhZeeQD9R+sQxes3v1HwPSZWuho2xXW+mrVdc01FtwEREaytNNwYJ0o
0TJakQbyybtEcyRNpBumc+mdeccKIGsYLjiMVJ6ERz2r4083vtFSqQbYZyYCAU2Vi3QuDKlpwfEm
rXdmrfxpMaVaW0VE4i8K+TZ2Dbyh8ikOEe6ZQattnHrK0fCrecy5kogGV4QsIT+Y6QVXD/eIdDO7
Ae2PXb5X7Rf4/ApLdpaKDyBk+JgQU+2Rv7sYd9i7pxcKzJizM86H/uKOo/FD+Npgon4CYwkUXTc8
omFqSAXaINh/6+3e5mb6AnFQDWGsNveGS0zyN77sgt3fYqKJLnAQMjLuTHTrZ5wC0FLpqNAFW7QC
M2455LjqZGbPanguHkl6W2jnybN9e4XtExtzRXSg6ZXCUe1upEtnxAQEIMBXzH8praUIDN5wkjWX
SDC/++NJxYdO62juJuMzSTNgYJTgjRfAafOCo1o6RQkSuPqExfEOJPJ+tjB+yGj8N6TtdckMERFK
BJHAih5DHnz7fa9Zu6yodynEy5M+WqcPM75pzXPUjYq8u89p1grbsV9WTgIThpF7lbSW9pRVvtiw
GtEgrDUrTHHrpRykp6pHZCpWSqaH1NlxePYAP6eA3CYJD+5EfEWg9ckjLN2ZWlyNTj7duPh0Nv+j
0c2PWRtEakiPCpBcqd2bkXz4VgexFvm4JaXzO3yTXHRZNCSCcQCdcQsUJkhTKBkvW+oqhE6uBpZA
thJQpXIlJ5ilviFVmXYJskvpJgjqePIpqIHJ9o7qVNoFKMOTvNI5FmaJWjqezXgQDkXqq/JFnaJC
A+2tkqlYhUEHDXizbAFN9s+uoxLw8J5nY0hzT/f/wi/hb0e6nzzzL+2OhX6jjizN1k3mlE7KfeeN
IGK1UzavSVTMRCsSA0ON/h0D/uy5sHNZwx7xAjNkN7Y1bvCAIfci52nbYCG8vqFOusV2lq8uBoBW
k7hX+0j+tiYstzLUUUN6Uh8ptxzQIr7jbxtwo4B1OW6caBDNMLp4JUsuaS16yKf2eWWnjFTQchM8
wxTp5cv7dkkEMwjuwfyGiH2EG1PBMaB+oluI3bk16QaFYUu6xOGI05DrhbxgdNeeBEkpAWT8B5CJ
3ZxLmGcGSevkwpgWy77nqJtodr63jMasMpQDVKq5RXOHcxhMZua+FelYBpR2yb2Osz1ojJVuIarS
mGgzcpVJLLsdv7iQeB4ltubjtz/o4/W/Eh+ZOAA4BW63IFlTeJSpYQXJBp+CxPbUrnTdYCNdERtk
c3CKRg/WykqTJYva8uF9RDECvugunYPCjvrM7S6lePTI8jPXL5GqxQV6Ww6ojfDfWZIACTSrfOL3
RPoQg9OaV12CP8oINwVzgoCr2lBoEM5Z/7RfqBAvEIomDhSys1cl0ASxiPbbYfzTjK4bEdgCuOWD
yYlmfqB4iFhVSwuZH2MdDYDcf7N16W/6wKez1VOVSwBL//khXdJPco2E3cvJtvgeqbkaX+YYl+V6
P+DOnlyPcsgJD7PdlTL0vz1DRvb5JDYTLau78id0B5YzyjdmQaLXoERAfPfV/pbNGcIpx6zkyEDJ
sIPY1/Hjb+UY29Yd+mcRx2tRtNQn+2h7pXFQc/tGjrBoV4ljsJkIt1As3WL9uLn7b7mYvEoxspji
Ol2QYCXBBcw08HTOZPkcfphIHFaHtRzX5bN0TTj95IP5f/dIsJSLL8XWTiF8lrC6w84LP1vz5wW7
o0ajrNPQj/3wVYNmmfF1bA5DfT4yLrEe3bPksFBvmn2r8fGgfvly65VPnm3y7yEvMvivbivVKVk9
MZiMZojzNBinPFkkeI6wyi6HvhXvPStwUHHhxzcmdEOYuZm8C+OyVkq/uoAkyjgXotvBpwJPJiQW
melPFqsTheyNouWOtptV8pQNsitYV5RvFCUS7q84IdRTUfkreWDR8DF6G9ohGmnc/YGt1e6wTjGu
nL3AD0tYMbW830xuwvsBQRM/TJp1Gp9q2ki0zfHxuLoy01vA3jPK++eSJw9tBSxmSFP1ML8l4W3T
XqRb+CbAK17/z1hzysI/3pNjQv5Q3b2VZBrsC37qftDwm1l1onPwG+/7enRSJxn/fAKOB9i795Fu
epGLqnF2xv2Z3tHW6UPOSIfHD/7axtyoz4Il3d9bdiEDNvD8MbUTg/bPv6xLQz5SLoiyvQoZwLbq
PPV/UQDOKUgjrukZSG1y8noVCY24LP9ztvG1yzNjeaRbX2T/VWdjxHKuayWZBTV1BsMI76hx6N3M
oY12u18oCZdY1Kv1gkVrZSZct90rrtMgdmWL0hluzp/lS2nXwogIdXdujsBU8KZM2IE/A4qj84VM
lprlBrzzo34lRPV61y6KUnEK1nuNFl/sV9msWgkBqa2YyMo0jthkQKWjy8rPtF7aZwiJU/L2jpTV
M1y0rxtzEJUMXlH7fvyfwwjnhDqHZPy8Z8cQ4gZUWNoFT6Vrh2Fc28XrjnBfiWsmtK+VDnU3nNjk
hcR/X4KEQ9+6eNCEQbEETPfucZefr8vveo5qDru63bVrqjXheulAfNiVAQ+h7eI1Eu4lQI3qjKjn
j0hCIXt+yiFVX9+sOh59bxQszPydn4X9soSl7HYPGFakJfWxPqKOMgToNsQHGo5N5z+WPLH4vxGr
JMnxEL2+7nlasqH6nptIHlHSMYdbGy2CdpcEexvf1rSuh9Mi8NAglg3K5+GUo9s2diCfKla6SEw6
jhWtSjA75H+VggMp3ZYHIU/fe7YDIwm44ZivH4OdTmG6vDkAyEK+Muz7l2jRelf4TZ897RTkdSxo
JfVJVtFUtzlZ9NLw9xIgJgSSUq3UobMJFTBZsB9QW11SyfUeqDIzaYacPeWg/7U20RcvQ4P61MNP
wyAT//2P/qDMmHiyLMN4VFqodfgfnr73/7p7y8EZoaTXWcb3TnDZwvazhYolyvYW3sIJseM069LZ
wtH9qB96J8Vjpl+3fLtdvfMJZS/r8V8fSVL66WmTtwWxQ17MoIKUgVSjzZsoY/64jQOzj3WpzJao
68v0Gxd1rHkJLedgmVxtJaTMm2eJTKEOFJ6CYREM1tCMx4I9srFBweGSQO7lIfmxn27GveZFdLqS
Yi5pKOAGo8jkJLygKeiCHbXwXWtXfevb2lYny0+2z9cBshkVa+SHH8eKn2hA4qkE3Ln50tAR02MK
yZYrogZmb9kV1a4cpCximLFhTFVP5LmjaFJ3ocdu4Z8NXxZojF1zlq7stZBCZwvju0rDb/VAA4UD
sdbCWr9X5vBbnYob2kY9sasxtz8QsFaQN6NqiAL0zd7GDPW9wOMeMwV9in1cP4RYwP46yR2cTW4G
LVvOvnz5GnliguF+4qmvk31AY1la0ao3Py14uP6UDIPQ9YQFDiYSzQ231CK3Hmuhk85PM6WSBNMj
Vc1w8CRC2Yh3zj1uRNB4pxQN/ce59rWgbmSUM4tGDWNaNg4cruB2vQPaNQrZbD+nxHEVsimb04HM
2Br017O4RBE4Fx1BtEs5Q+nbCcPdMRj12dUI+skBkqXbYdxIVHy7PFMKqXqEjGrf+z3+1ioH3vsb
f3PF74+sehoJlI2aVc3HpMiS89xC9I9nMhIvgtFKRGpK/ZUF1Y11V4DWJylc4RyU8Zb/+oxWHn+k
azgHk4y+vRirLatt9qHXfR3JkH1opdve3gKIUg6v6sWAAwo/IKIOBlwH+1/BnT3hj7x649iwG0R/
NMXNathfRs0yoh8miHxfEGFmv/r0tGSFlyh3D/Pyu0BAIcVwJHXTlyLuioQpqipdT1mxs1OZUItL
dAb+jaRXuZhGuHYQ77nr3PKZGwHfRVd01/Y5teiMcVnkoSPKeGH/mTaGQ15eXlbr7hEQz71ZokWH
cbYBY5TmiwtDzgtCgtdCB30LLa/CTvani9d14SGmaC3hfBx3nOq5SQPB/uSMxLXLRNwVO4auBVTz
aYsYGXsJsQrQAm8vCZo94v0Lda96zSBY5l6MjRBBm3HTiwqfFt9L6KP5LS5GpV0PjwkEiRhhHUtA
2r2zvlX3Ym/beObUV8omMNS9XqDkQ0l2RaHSm2VoC2iGDzKBeUkqnO+onwkpykHs8yuNxlhXreCO
joJsYH7Pou84cIwXAH3ghjTc0H8NJdddc7P4/IEDhVVpP3cZUyiUCHLotxqZ34HF22jwNBfIPp74
2HKUQBXmPxRDmLHsLcDvEIyWNgQ4W6LMlxMrgxJ2+9+Yz1Xa/Ar9P0UsOwEJDt9uTHmvLR/1vELQ
fCqGdN9SP/eiiSv4gA++JQBH7/HJJbkZiZgpnNuqZ7B4OVtHMA4T6ylO8ume7hRbclEyAy6mW+UT
lNYiCQAUMZy28K8aMWhcPs3lTo4xxMcUPMQdn1Pj713jS3ZdX3Vk8VA8n1UngmzJDenN4X+DJfQj
aERRX2vsyqxIm9OaTZuiRCdViFtuXtqH8mnoM9U6tPjpQrn50WLvWNOkT8poqPi8B0B4QEIpOLhb
kWzyBuGXM1XOLVmY5d1oOKfCTUVwjpLQcGHgDMleZRxGJUbt/k4ZFh+c+1JrGMpnI2gEU2oKavyZ
5PyFul7J3bgjx5ISZyYxya81bbYxFCDR2JkTORFemlTmX4Qx5NXq0A9ZsmiD4+Q46wr+iZj6V53i
RsMiY+drJGTFcQnPIRS7m4wID8AS0Ivz6agO2oFg0Gx18YQzhrCOXzA2j34A9oeghyJ29RCVdeeQ
Y7NO5LCrQTbqEXbjCE348FW/AqwjbMfKBoVZVGEq6wduncbtfTP09Ee1XCPNx1UC061n4wPfs0Yx
/MAmsD+6UYHOHljB2e+W+Br6g7V3EP0wFlOa6kIMRqsiy9DSCMNsagdKHVEMdqfBXytZg6s95Jgw
1Erw5/ewyo30TE508kB1UMf6Z8e+x5KecHYdbmN1afGsqDF6/2cUna3qi6WAhzZoN7mqn2M+Cd+S
Amsz76xyQNMKKaFopdMrHrtRkUWrlBUyJEvS2TnLIcfij05vhZVTXfyWEAFnof0AJ755LsAvbtmW
kgJf1YDZN8ZbTsqZYta2alIKOa0nzGqfSufED5ZnfgAU8I/3ZqbbjO/6ShXuLQutp6a3i6tjSpMc
Z7GWqi6fdiyGsElWEgH70IOSKetc045nl7GRH8zPIDm72PLSSf/W0FRizVqekc74l8EUDeCRxjHP
BlXYqz34omS8wUGwCESJZyzxkoizpy4R3suriXWnkIqffANAkFVnwx6mFu3lZ1quSFOYEtk5VG6n
HfXsxI0gteScVfaDwPacEH/4hV9T8bbMkHDTwBCCwFUqJpjGJBN4JzyWOM8jwKucH04ON6yzXDbw
5HXKzygZaJXQEtoWggT5iAKMKPbQYYxAUNkbTolT0KYB4fc3ErQBFHRwm8juh8oZZOt9bSzFScvy
l34aO3LX/neHzYJPlWinS5VeoacSdH60Sy0+/QYQhDW7A0YVPfaKmblAknOTi5g62uFEYyZT4mSV
HFObmyZJ8cwLo2P0grEMAQ/pcn37GTF/mExhDn/NgjU6ilZeL6mwvRbeg7E3cJyCFw+TPjYsyos7
lvzQnWXzRpONv06efVlGn6+MznFPYxjokS7VLIaEeRnAU9QYZ8y9WPDVug0Hm8KGjkI0E8rIrKKo
43g/BNbmihMCjG4U0QLpomS86p+b7BdtxicWrJYuKUvg2ucV/Xu6zlbajt/5keRr/RO3hi+Oc8je
t38QBvMLR57ACKIjtcre6QXW87lK/KtxIznDwxROdD+y9W1I3skx3i8mH9DHYG2NThb/t7K0htaR
nUIUbd/vWZcjBdi6J6mrxVU0J4/7ESwXsN48PiTK0phIzbTjDtBIF55dxVH6PkBTeSDnpg2shpzM
P8MgY+HDaq3drEntbK69h9NbNffdKC2os3arB+DWW61/jdn3BQ/j3m+H7A345Zi7Em0nqikd0cSD
OwcLwn2VDrFp9o3dmg/HK02J2++3RKbSfC0qqcoJsPr9/4wFPjJ+1fVPQYDowrfDRNtcfyFZWijx
81pW34F0Co8KKpJ1WEYOLolyMbHxnAXilsfA2VxwOlSDr0T7BSlX6w3GuDSmbQ+LpqFkS7cjkd/w
0tzjAIGliaHvJ2rNg7gjfSlduHDTw3qhzlOjcmry0rfl/SZEkT5LOu8MXJWqgpTUwImJZfDJ4LoA
nlf9iCAow0EPYqSv2zynwq4+IWEKRoCi/6FboQHWtbvk7IX/lwSul47c1yLyDuOXTTfV5nQia48A
FWJYZA7PwXO9KrDWD3in+obteQPI+bqomP1dhQghPfAutISbYe33WOcCAEYm28SthGxG5ch7MidQ
10C2fTpd+Z64V2vYd+lgdfeJczewV5Mj/jeJ3porPn/3Yf6A4g/GWDQQ3JuZ0Sesxis+2T1Nz8Yq
tWlGIh/c4zFY8If+cNUpui7Ly0RukWjUhAD+Xf6yAQUkVKxw+3L5MNf0Yc60Eq3JJD2afypwiXlJ
RPmTGlAvgEyjail1oSID5Y6lpbRC/lkGExeSgQZK1vupt8G285uQuG2KkSVJIZRYRPK0z+UHAYJS
ZJrgvvoELyRrZuSCK8p5inOV+yTERUmsOOmMm2yVLXn9NxP14amheALCnXMZQ5U6FW4O+7zkmAGv
2MBGjl57QeZdfpyR8VLbxk+w+Bx/4W3lGFWVIurfwa6TvF7HPUTFubrrjQoNAc0yhoGywa96hjE+
aa8kKVRwdqKFYT4l4JNB4tALbeFJqUUUFQ5P9K1kLp7MTJOKb2t/knAcnz/VegRUwPSQW17Qjbv+
Ch4Xf0v+uR1nZsVNzzKCyHj3SivLob8utkeuIE4il+TtV7R8YCr6627ZAC5hRjsHmsJAQw4TiQbg
nq/LNZS4xL0akPLu69wXPO2lJigbk8RwpTtBXNqFHpRMF9c+I7r9vsxSfbA0huB+A0PCg6vAwl/z
UTtVLsJ8Ne5zVqPpVOGsgo79HCGpYMQ2YhXWbII1mbn6HSMi2rbi0DzzJqOFMK6p1zLEua0AeuKS
HRnCtCSYWI19mGNHyO2DBOqM9vR9we/1WXSB9OfneYhwZOYE3J07ynYE6XR5xePFEqDtW6aaFCDt
v/4Xl8L+Ick+dFqWqnv91hZ7DIFVk/LEiINb0UpoK6DYzwc3dp4My4pEZnqmEoxbT1LGHMT4VdV4
SBiAdvO4vaDywDyfYn2ffeAkeZUtDHJ9jDVulIhYK4v+YTBinhr1t9YKW8xDcvXLdfesGK1W4tlA
eZoZ3S01bNR2fCAq3/onGA8uKng8W0o90m6SZOm8WKrW4mbwLqiu/Iv8bCZ2H7Ke8+uSWnrexvLR
RNS6clG9PH3VCXLltFdTeZ0Lt3/7DdQ/nZAv+k5J9STV5Ii4zc0ynihQ+miIrwpulfDy1Y2xapkG
ZXrFVxpSo8aA7ma3EtCXr0EeS/kFD28Ucif0GfLS3h8BSNE4FYJMzPx5cYIjbt0gWbeIPYOaZR8m
op6DAWl/YT/kU0/5rz7JwiZOheAifHFmWTjkG0Enpfc9fQMJQ/0YAgOx/dKsB1/AMEKKukJqllda
dXWL6y44+JADayTi7AT7TCO5bmMzEMKrZIehQBEu5WKrrk5ZK3TOe8qrSnfBTrAvGv+k5FNCLV+n
a/x2bNIkQutRGx6ealVI/Y3lIgWUUKPXQucl/44zyJZlHRBthLDPxfF0aGnJhlISq2VGuawELSoZ
MZR3VJjuE6uUuzVgZxUez9xiAYtPjrk19PFOnuxSHuV02I7G7XGH38AnkW2sMHd3JYDpsWFrfOPe
XXT9Gj/7CMc83ugEtBESgFctMiTFr+mxR0TaH15rR2o3OfmyMlYRdVPQAqlmswRk0j9oDEZ6boc6
zzgn7HlnjyB/nI69yzjYdekTrcUbs8FUD2Kd5HE0niMfaYGx1Lkmu4BSFda1JIa8QL7IomSJFjyL
Az06BmGXFvStUehCEoB8TvgEa8WL9pLX8EKXENWjLYFw0EBkzTicG7FibPpiUbSV7P+/XHPHmuCJ
RpbWTcngvgxk92r7IBUR2iCiLlSjsdhVkPugqgNGbfLRck4gi+x4xvD8pM2fnAZrU352GtDfzTPR
WlSz60Sxf8bj4HY/jVseMNfDlp8/GyEKNi1ZATVRdq61hl9oA7j01TDVfwihjId42iIFusOthQ3m
uMswYXMZUaP840RFqt9K6uR++GMG7Xj1T+fBA7lNDa5mzPjpMs0Tu9rjzriZOi3jiP3+fXRYmfNg
PUiDEPK2blkoXoaDRyR72jklUvTEOqiD80VaaPrFxJJApgh48PRzYpzKyBySRVgIIEqL+z6T1mj9
fE1ikDDx4kunwxtWSv/OvAVN96NqVgzt1gIJhyI/HPCbwRHsgYRpdm0z9cxEWngzXSPzrmQ2sRUg
+JxvTCRwN748dvrbX/1gkdh/4DEIfTo6lbd992fW5i6htJ4BUe3qwgQ6GDpNk9CxjUjsE7S8ijKl
LP1vrvAVrs/EM+rR9LYdZsXlF2MW12SOlA/hQs5edFCGzHGY5djbTM5CGtj/dETkj4es6VpFwpHA
Nx5nGp24LAuaDwOR5UJJ3mN8xdfdSbqFYDsJyXhj2kw4u/pYQkLAaqpIrXoFIYH5ZULJNBDIRlUw
g0QViUq4RDtHSAIg3PeAdgVj7xO9NFN3afEx82zEPkY9swQePssgdNhzGRCOoPaWmDHZLbX/FFXi
q663/ULDQWP1SJSgL7JHwtGnbKJgu6lmfV//3uhp5ztgVA4ksg5PHai98oRABEIh0CvGKT05xzMf
hVhWYbaR8mt8V9f2WcgDLhIVo0pby+eMoTDWG2UiamH6wU8PzrB7xn16hC2GkGGKU5dzo0E7eslh
p+5+fgKuf0FFtpltCpI6qYscZYG8DtySn0j9UKWo7NRZ+ytbXxBCanxmZIvE360FM7E/P+wuHVES
eKxztddPhU27Td5T1JZ5H9wStf34nw67x0ph1t7N9Qh7Z/rCULNhfjTKCnXsSUXJup1R3m1XGq73
CQnNEd5WDam4YJaCFcl2yHi0vzoIai6cKz+fib6+wogRISH/ZjNN7PfmQevZ/wg92PAwngE4BZHP
Zb4nVCanxuFc4ax7CS8xAkyTvl4ZFQvOAoXDZQu/6osjKvkgSVrkKbN/CSurDGtkne/DeBPA7Ga8
OWZq7NWXeqWvPtQayqvS1DsFq6J0jgFVAZagiKsF+1RfID5ClS7gI/DTuY2jDWFS7GxBR3xr+aH2
koYP/H+pErGG4f2Huv0+ia18BiaRIGnjEIo86XDFk/JG3trvNkDRaFhvPG58Lk594wuWwDjQ/sfS
S6RuaRqPXo8pbKLdZCsXV3ldAmNcJ82h7Lvv6F4doBfGgJPp1YC4NXu/bVPa5XSJFoL+2vjeIVJn
OJBn+iKFfcd3RxPZ6TyuST/AOKJrqazy6irApMlTpI5vUqQ6MCgdl5I3fVCndp9huqVdwCcLL5ty
+yWPNOgob5DPzZKgIZCBFI0sONOm5Mx9+r87eg6RY2BZzpIuxMFPng4CZzb1bMLFzy1XAD4VENU0
A2gMQOVJwgiMbSMqIOWFTd6w1CFI11IhzqLvO8UNwJXrOem7UxHcs4/ouzgCSpKNlv/ec+wlG3tc
hKSKn6N+6cuQj0ntywhMpEpxusyjpAEL7+2Lv+kjzYMuXT9m384Hld8xMlTvH2+VeYVKtK+JSMa+
zFAh2BExs2L78o9VutSikT2qItXpkYORCVjxeF9EtjYVhukL41IKgmFTh6yI2mcC8Id6nKJtvVle
TRIjr2kWu062pnNceejx5gPxoO0t+Q2KPc7D+UPt7LZqpYiN/x8zMWToiiiJoi2c6JK8mOp0bEFy
1alVqUURR4ZcWMS3NVPyQ37pDjzUhYcOlRiYaermpdvL9JLnYckpjvPk+6gY/RIfzVudingDZT7H
+yfwFccsuBYCi6UAwatwEff2kZS/WR+QDY8Jw0QmaNBt6rb/aeF2ReTyZTKjDG3IdCW4dyffAGg8
5KWnOmoLUWmIuhQrkQo7L+HZnZorl0PTxGtxWQtdeEeTmtSy35t/llc9fCrlJ2XdU8pAxHvLAs89
/Ns9lSFY56+phmEfr2iW6FriLJ4R/u4l3j56jAQG6+gcgObEZStsDs4korG4FCADS1YLPCv6uls5
SAwocSsF3PSXpBYXSdgJ+2EBg/5kzSQ5ylnMjNqdAvIV1BSHDnLR6CuQ2+PcKFYXC23e1omSWqf5
NISt1RulYSkdHnBsNNC9bqKXIbwNYo5h1PTN9+xetDgjL5NEniFiEa9GscL96rjfmv0mxXciQnIA
8p7OThgjTrnpjKVZHv4hjqqiXBIR6tF5hL22bPo583mTEB37jXCJv0qX4cTNz2EW6F0Tt+Gjk8sQ
+9Bls3L8jvP/3BYDLIPAVHxTOYT5jTceZjpTdpX2SSyNfRZ7XmPOFBuDAiDh6fciBw2pmP/ojQWw
++b11F5ANt7wTSkc5mfRyUDqFLCwYLURTYz39syp7LNLXhVNaWTAbKTRNwMTggIyXLzEWWJ3EM82
nhMNdoi8DNVLwipu+PffFX1n1dAcqUvAlTzgDe5uPJz0iJ5IcZeX8YXDujBPmccct8iXiyS53k2F
MMnVnuPiqhBHMjx07efzu+lNj8tB4TSvRdi2rOd7sFVZ+HndHKnkHLeFbLmeDdPoZfvOUOkZ8mHR
XH6CBK9P9VQG7QYPQHLuGUsWKoVmEPPVKx66vy3sNbsbVIbrmpQgaf930wZ4Iely4dywa9hIZ638
qhKIakFf+5zNbttyu7ASXBjjaRkfUVGEKYqcnIgv6aV1qnH0KX1Wp+5MBezs/sVBkIAVuSYhUPFi
2VtPsRVjvgFp73zjHbsAH3mvYh4aPUoZzTQZzC3Jk78RkV32E1/yLmZlzK6tFJt0qRJXF+esWQW8
zA9Epj8L7bRN6sKaCjC0tOsKv71eh8tFuzSx5RZ2OR5C1shOi7Fthg7IvoX36AhFcSIPsTiaorrz
autwgnoxP6V98hwSm+ve5Xm9Oqe5pOIwyFatBopBHfHsUaQghoKlAPTYtEhFs6sqcDu1tVbrMLrF
H2fLjtl9r4xnR2KkF5Prk23NmmdXJAl2su/EzpxhlFB8RQ/mamlgWsKhOMGdosn8NZT1oblgm4um
jMFSWik3DsELmD/otMIeyflgBiNqhPf5is2rZZ6FN50I9Q5RwOZ104xn5AHI9/UBbZgxfEhGJ90Q
cHnaBtS8Cl6qh6GtAdY+XZ2speLIlMw2v13xTNDxLXWqtcp4hhwyAimGN7C4nS5KeM/Y+0vmDcx1
129E8hoNUU5SjZ76hlSTV+Klj739vvbG2XnxuIuXkEbOHLcq4aAgML2khEyFnNXPCwypDCCmQdIn
i247xxMjQIXNQxwy+6MMUFXlu8VuWL5rfSfnkkyCzk7hiWE4qf2dXxn/bMg/lQaXsvaNSEuCKyU9
oAnEHTM9wprtqdrMH4oAaq/kD3EaFVT/3oH3n5r3M3maXrH3A90f2IMYSgvrsC6bJKHaZFBWyQ72
yGhabJtvBrOkrDh31mtSsxrgOq7vo2CSP9RpDpr0nZpAAfh381PE65v1MJOVC6lOlOcLtcqHfzdh
2D5p4uPve+Kym+elqWZfoXzH5IU41EPYe0LfDdEg8PxlpbLbJ/2ZeAukjWmy36UzAKjyhYPLyYdh
8n/6EIca1X9NZmT9/JLrEiO4p07sVQzzdWQc1acGx27+uQnoPQOUn3joIk2JboLC+Ngm0p2dohtb
8GVkBrSzYa56PmUFHvnmCldEzG7ZhSRKJgliVRei/gF+wLCrC/np86HGghvxFsqamu4AvG9A+lRR
XB52HbtGSx9DmP1t194CvOg8GAyt7en5MXMu5iTwZlWwTaVRGSwLp8F41Eu/kAJN1pnxe0m/vA6c
X0ETQocCbtC1rf1dpnzfSAAIDuEjYmQ7H232KpKytFVjIKdg3bhHrSSRSHjAEAO/1NuxSd0gJPnK
pog4z4CSqSUBo4yEJlcE1Q+YjtrlPqQllxsFtRcSl0jQKkvqA+tO0IB0ipcTWDYqL1JyvV15F+Xw
zJmXKipznYlzVSww5FiArqDqABymzOalRuhSo3rxGh1P854LT40Vav+zkaIfg++Kz8Jlo/m7bkML
HCP7eYAxalF4kHqzz5RlSCadzbDVd01Uo/onVFBroXnh84J8AttAGhWCOg1WcbCqTwR2L0MA3r6B
HI7Qi+jA2/uUDg/I1zZAPGdxapU7AqMj38lK39/fb3lyuby05MkZ4ZOBuV62pPoJnhDlRTqHA9pa
995mk+fL4TprIPEq5vuUHngQ8WrWkVl3GoBTcDhB5YJQBlL2m+XN1VxlB5kN2sRcU+avYggdctrg
mgOYIY7hhFdM3UHHeYKSOslLbUadAP/fbD8U6Q4smrrbUaSUqveMwPJKRVjqk5sQxRdS+3E7UBl2
ifj7LzjwkLlio7XP+CHEILuOnYZUPJYJfz8+Fyr4ja7OM4CZh1ph565CtbJ7xsvmIe2k8bRuqQWn
p0W6YVW27hlWe7ckgveKXkZeRtDDVVn+eEuHq8C7WbT5ZpHie1FsfGF4rWZLhGmw9tAxudD3l7vM
adgK2vgAb98g4GNAoWG8wfGG0Zd0CBtCrqpt8P4zLFF7VH+HRU4YuuGNqFCbO77pkqWhUx53FYSi
G8LcgTDzobrkOOWLJZeWFOrPEGtRTxRWZ5E7KOZTdO/0R89VxlifhGvA+XMviTP3Bq6kGcj5vaIz
WObUHAUBTZxeCKK2D9oMjWVSFSi8nCnZ4DdlzEbrQEp44uzVDc3K5JInTcTASKJelw0rPv2eO92S
w4rWO0R4KoR4hKvWtjz3TbxT5eWQ32uNlf5mKXcHEDFKnRDhByT1VGVJfKtyfKUk4StyWPOgtQf6
zbeecFz6U6vv2NmQKMrcFe6ZtmZ2X+zOrOiFuJPy6gZX1Z+U9pdZBlYyusMp5dFgpeD+YGqx/aV6
+YUdstIXoFhhgeRj4YcB/rhWtNdkuvkJQ9o8CA/LSoWzi9EbmAnhEze0pIfWWickHA65xQko8JvN
hdZ3w01DceKbkjUQ6Ic5jyBCi2o5LwI3/PGs0sEERAmmgsUri3amXUrU20ew3IiLa/kGfPCvSlib
cNxumm1rcECmoaM+8NvMdgPfVAORWF2BAlDvCNHGkBnJQv04N55Lg8fe9Wkpczd5/l27Stc3Qo+h
qi4nmB4RWIGnk+8mKuReLJ3il1LVt4/csackzlLFUdJVVoTPvFX0qlu5NgGPa4c17njJYaKLRBn+
KvFfk3qDwiZbMPBZGhricpypDHPAC6Vym4AyWg3ii5wqTWhlfSnKAHMXdZZdH790SLJ9vUAo9NIG
2RiTC23icC4/xI4PD5O2zR+Ldwo17WO6ZDDU2ctxXib7oUkSabqzy1yQIbkTBJ9NfylWHqKMUliv
RW+cSHk3Dd6Ky60IsJHi0Wcj/TFXWSWATGMl3OWs9VFI6tBqGWk4KLmP2gdPrjgkpUFqfTJPU4Ss
mAdMpjCsE7JMb7IQymmsdiCIyZVqxiqgfAbhUySIyg4VGCjOntuSWS3V1aiEI6c/PxdohiYtUxp3
Vz+/mdmJylbl/m4+NjL4eGIqNFUxcdM1se1PwsBK/oIAPyyHxoudJIYFZy2gJ9qFTczmrUsS8NDN
XS6qjyLoj4gpEuhuR3y+5yCAsYf5/4dVxBacznJYSgRbPA5JVUeR2DycAZcIrbCWP6x3FPLA0huz
jhOuVu3QuDk//Vno2dKIqvNoPUhLSvQb4nIrc4GkKYfH3B3bHobmL6WTaoHbcnCi3h2UQEXzHgYd
BYJr9lkoWpRYtEDNN8Y/TmyAKRHKcQrz2910s6KhAxIebI3IQ1alhlNcz6OT5aI/I9r1aQkBNvCF
/ugj35dICbz3sxijGv280/5fE19GyXma0Yvf/yFoep06zpPOzr+DHmi0EmjZdGTvHtbKbRTUUpiy
l2PyYffJXnRUKfNPTaDKgGrTivTjWhlYTzzpi8cC3HWRF1IpGZVjvR/4EBTddPZmoQCLxjh29cfc
js6gHJE6M6Il9oUBDNRNdPm6XmYvHAncdJanOawz+hiitmKTN9PKjA9NGwD7ZjlTnO2zfvEeOVpo
8ZGdG6WNYjoDrZRuS1SVyZ4l9jBk8KJk+ZMDZE3L9uVrt8SeWBJPKMv4733kixX5ZycK4IVtHlFL
ttN7pZrADCU3qW63I7USjq5hlqzNlaqpI2hubtv+Xi8Wmq5qVQ4YR0pGBeDHI+F0UIvhH/1xl95H
BRPZJlUKkWuhdaDw9kjNLsl/foDTkhEV0ypfEQi6CEN98XcqzAqgMRcLPxiQIB9xTDZtzSDkEetJ
t9JrL9AbuouFRxmtxtOIYS4E3AQAziXI4AVf4nCWPAzUIK6FgpIjID9d3iZeBwfVmDIC7mlcyV9I
xNqC8UNRqm3kATgfPcwvOlp/9k1cKHStp7JdDF6nHAwzbc+VDpZKnn7l6j3AlFHnEz02rVKLr0nX
h9w4jJbTOvh5EQ6jl5lmAE4vq2T6NtGC61iGGw5B/e9hec+UXe0ME6CpB7NPxMJJz+LmpkXC+KSp
pQeA2mSlmXZddO4FvFVwjs0CsUkNEKcrXX1ce8bj2xiSjCN5OyVqYqU1pF9nnfv7l11/LiCLSl+o
cAU8RDS3pUDczij321YOSGJEoiwPMOb5C3PzGwIoZTR4ZQridEFiSrpeISpvIgHJ1XBKPl+FIfVf
559aby7rbVooOR4bvQcCWWpamvU4QQ3JNiF0+sAtUBE+wVZUzb6VdPhBPapZSX/W4nY4INXBRjrr
tMB0ZvC9pPf8oV9kg8MhIgrrsk7vQ6ctthDSjS2FXNrxu4mZIflCSJgCpmsj6nkMAo+eZOwTtENP
baLUzUDx68za84HjQm1dBU5lGVOAtEEppuapKWqzZnHyXCkRZ9pzhXx7o/+PJfa6nvsSNbxnIoB9
zxrtcsSZWgRpbRQJx7rc+LF1I2GeVmbAeSs6LCi98Dpf/mGvboop2JcQ02i1GAwl8sT6ci4PrLyo
vFSkG15JIMu1Vm9/mazjRPlLkKZFl8BZ1nD2pNwveLKHI0cLyvP3SIwhV++YjGJ7CSLzeYI9G3eb
kJEYH/NhSFL5aPBW+i8TmMuE7fReAY+cQwzlTCfrjRU45Fz8gqIYlvXyqHvhY2m2xwewiMinmqQg
595axG/GWdJS1zdIFi/Kv6YcrWEIpPlhqRjM6MmKjpy03hpCnuy0T+dKQ1rXNq7rMWSxFDh5J/Rp
d7F+jgYvSIU2I0y7wASrV6DlWgoNKg1u7ROkOiK/35zLIQ5imolTii+Y93XjMEY2kzFNMVkn8ixl
rG2k7ivgb8rdxgeMb1MpCnYlJYo2GwjSGotP8pZJ4Wa/Sw3GSBydmcuLjS0pLmDuO4I8pFDDnUOE
H8dY+cHPDxziKLMPm8WFyFLMnsbByXje2nm81gy9IdT8fPMbJJTyMoKRwQCt2nKvvKVTtgVS3uq6
CZ5SfkgEk86ZGTp3nRHi8ASM5XUN4CtEpyZT37Xc/kQPM0qZ5myHzuuVDFmfRukBSOtNMaX5XqHS
vJq5gikTnFt3c6XLWu3pStq3Y609J/M7jBAi0a7bbOJE1yyBqeYdzA4/HbzfTNsfn8MM8Ol5+sMS
Q29WlZApdslJpO0n7G1aesBhciJjLH+aqLSm/wsAFkrBGN0KqNqqtNNnhpLV3JxHEzP02pSrV+gd
BdDl25kfLXGbZWI7jYhtZXcLyOSgBk1qX6kDCICmrYfW7kxpK6dH9tJ7O4CoQhE6R45ItV3/sO3x
fEoHN6a0bWHoQ/40bhpkiNNVBb5LU3yKRRUKlpxQvdrNNmH3qjE7Kj+h7kEHejh8teA47j9YX/yZ
//tqKJUVrreyBMOe2c0A2eHhM/ccozldo3sw36Bo78qHRmuteQsZbfaVXrzEgTJmelgRbIQnveb9
g0FUw9FaYZGir2TAbliEX0mtCtITqkeL5g62dB8atBKPibfOvv+u6GwWYJajAErzNmmZ2/w5nci5
x4uDOqSDYTJYUAA+kzbI5FBkfhNQCqNNpgSLfcN3GPFRnOrJVHEiVgax4aGAYI51A6hU8GHBpBVC
neYpMf0Krit4xlJ/jTTgwUIl/iIKMoZNgIvo71ECv/t/BL2dFzYJsT1zr0N3Wp1wm0QPa2yc8xD2
l7ZFofpPQsiuxKN5LGtCVuCMkAfkzyWMMoMM1hmrpVcFGsZvEz8RGJtOvXX8MBTmk+mIll4tMpXY
wToT1F5AQp1SbcFJJYGXMuvV9Jt8Zkf5On9ZrKKZIgEhkxMMkyuPLseAE2abrqkvHgpnq8VjJonM
sTidcs5XfLK/FhOkow/wf3V0NPDhs6SP9Gt1H91ODPztRBYaivKLkTgLZZHlllrxRnNU3fCPDahN
NCsFCux3CHBFScThXiqcUcvivn7m5MiRZ+33YtGHZq3WBTaa35Hj4D3rlL6/Xbd8ns8uQ0PqiF6F
fYyZe4NiokoUkk/Xca7dRc+vRpQa+CGTTz7dY85w1gEiJ/IydcE/tSa08LXuGJddbIGumoHtjqDQ
OimyvI2yBMdrH/t+ft1byNRcerSGybQOgFCu3MyyXDaCHToDiBYvAZz9kM46aAQuU33sZrjoex83
eHIr2Qrc+6Z07CdwWATTnAZJ2YQeohY4c9Qv1CrWb1pVKPIkJPvy27W6foq6aVi9YMKWa+H1HYWU
UUBYIghcddlB22HOJ1TaDVd/IIEDxYLv4/2m1yNruuWac0dt9fiTeeGvyKv3r1SmHa7WK/gcHRjj
sNTFdNd/RU7WS/nnMixc93OXEueULGernb4w/HrNaSYKdfmcPbRsg/7Nk1DhUV9soy5xoGbIIN1R
lO9fkwKWGoq0jVLhN9E9Z9PZO2bS6rkK5H7DXgVx0lmOHJquEzdHLnYzZ0gh8ce7gzLExADnTVDJ
nOFRAlQRESPA2icRcNxkm82MNa4NeioZO3m7GnX9FOYIHvDtoYkPGMRzRS4tNd4MF0HbnHD+vxDq
r0ukwB0wUyVoc2n+/OJaQOj77CH9IhzxVBCoj8fabJZkRi5LsI/dipc4cskZcmDd9pqha6/+Y/RK
9BUlIc6NR6HVCEGaDyfaV1JGet0qfmrCSBVlgl4gVOVViiCQXq+2MWIm4NN2RAFOdGn6Qg9JHVl4
3LnZJlWRDf91MvmTznZJVfKDB3aZPePbw8ikT7nP45Il6nsagmWvS/Nn8137irAg2pWXRq/gwaWw
ZKrQ+NMyfcJ8emLUlXGEY8dLNx1n3bcx6OxSYrkuwRz8ZMBN5j/wYFxIbuj4NjVH2caG7ffEkivx
167ebeObOepYQ2V+mfYcxR94mAhkN9rhfJG37uere6VM6pFpyXBjgA7R98EvxxbURK7Dm4TsrWc9
KGg2WS+YK/vHsP1RoG2IMuxtrq0rjPHr29sYh4C10Gs/WPVF3XOKYHYLRHgl56qk9HFgJRcRi9Nd
7LA0zEYS3+k4SzdI3VZyf807RiZDI4ksrsf019RUotuLQ15aDzymB7dKhzjEcjfpadTKUVcaXqne
t3jeftowPhoIOUhYBRJ//tpYoACU4dFm2cxNzjWkvXDi6If3NsI1ebubP95AC4kAQJazee2kqmfp
LyJxU3+koFJakLUOVCLSNri8Z5berpxajiQII/l/UoFBeCBQa8CisfBVLEl/3pRTaXw+RFFVvEXQ
4NAuwLQGMz/htSvu0RJppaFhmd9G13rzOME/TZzjhOvrYL7pJk1jDEco7o4GQ0gjV0sbwJeg2Gms
jp5jL0SQDldlabvit+HWdAqvbncCko2x6kuny+KHyMh+aZ2Upweh6xlEVzZKvdtfnCfxQCiVNMjy
qyhbrslT4BcQIcfMc3U8HvOmnxfIiPDB3JllkOAGFFcfr5y0HX9MmuLSp2FBdkZQSToS/UtKLT2M
BT8SYFtbJNIXdoz4Amrfb/8Me1Yt62P9QOiwy3ww3qVRqcoWWZD+AeivM6P1MyYqUcgQ6tEVSuxD
B9ZRBIZxOIVBtbqlC3Mbp9PUqx8E5twFqp1nDuPCJDugcOGD/m2HJLzPhogpQtY5i2pubQDtjYIV
g3aDFF0nQj9RfP5qS8vdJlDdBNi/KyJXnG4OT7nyZ66LZBe9b/wnmL8HUnMR4d0xx7+kl8B/HgFH
vSJke6bG4Dtcm//SbbPN81ngZCRul6Ve4iYS7Si5unHmAOblgxrPOj1Lbnq8eDNO0JgmIitI5DK9
FSFymLNpKay1O6p49ouzHqkJ4gm61VzLrUjXIHAyKvkndmCX30xt30ZeHL5+w+jLr4tw51kb2Z6B
xxNoMFeqsisy6KGn6t651XG8Mdg/4PMJnYdD585aH7r+k2134GE04KCfDjbVzvdAORvjcY/pu28V
6t6WZVJvKKOdZ+XreMPjT9R5dKNU+YVkOmaMA4nF30SyQd2tFjl33Jbk8mDCgJE1hucxBaReXJSS
0Lo29Hcr0QYr6O7Ta6Ory3DtrDTuoyrQGWZtYapm/M3yeIHRVjkPyzcPoxkKB2/nUGoegGwPF7iw
83rye01gZMW4BDKRovmLRnPDXakO02eqWxq5DlhOhVj1EB7bOi7eYlqhS6cXAemBZQYjgejXTgFp
ZgXrg9UNI4mYVI59xVYBd8MFQ43wtIXmY5ktw5wlmXMYvdCun4n+gGynO+PGw1YfJ7eIz2va8euN
J/GUNN8mvV8CAOeSjGtWxHx49CBswkqLf0zaMgG4jGRAJ59JvQyHJE8RrDXXRBtyKRmYcqlE9ivA
At07py6nnUuVbhqFZaWVp3jld1Icz7XIb2K+8JEPTaINXft0RixBGWKdw1wfD21BpkL3BnPVc0vq
DoT2HEYNHs90+AAjAgoxUbx9uE1Co1yOk3uzAFkxGg8d7Jh8vvinMFy/xSAdnfc3eu0iqjmg9QuR
n3X/EprtxD5gF+zHERR51OimdyFb0VCb5n/zH0iP79x+2175i/z09JLhGpIPQa+raSpQsKijfCQm
Jb9SZhDY/QE1zKig+BRWR1p+FNv7a36SI81WF0PSoWRwa1sfhi1G6B8q+y9Bun+cHJdj34VeMVHx
4+kO/rvdGilC42i8VuuFsy2jkso7mObWYT/63COtW2Y+0tgFEDn37P3aV+vmVVnDSewMbi8JfUqE
ezm++F1Y8cac7PR03clgOQTMADUMUhtHAmcZbvcMMAmBi0KtWKMbHprwHG+X/S9/ynlM7q1TogCb
BZVxArIvltRVr3iaC466thwUYTTxaEWOUq7jcXyb+THaDuN+SMGyTmEsQo1ufdOnysKXJzp8brg/
943jDvZOardpq3MTIludRCrJqvKnW9um8d5UwYT56Pg3m6xhv1O19Jvp/3p6MLlseH1IjmRr0kvP
eaPe82/Gausk0GoU3vRxMafoTXP+tPPP5ndPgZcbWnrFv84IdO0YKnFrh4e8nO8DM6m0k69p1/h8
1mOCqUWG1eImyViHNSzcWWXOlUorbe+VPLj7gjROXLFMEC96Ftg2QaxT1XetqsdNbMMD12W3qHXJ
NH7oKxNr6NDlDkp+xt3Vn9OV76aSivlkMs3JTUfLm/53iJxSKpAMLEK7YDg41eUlETO8gt1pHNn9
mtpEhD4BmXrxauCcGBUaFAzMvPSQDi7AsEbzKQM791VBSOGiDdDzjfECKjjqH0JTTVMy78w6qkeD
Ydd1Ktofq/OWM9d6uKybshqAA9/h9wWraPc8yqPQ7QJzCJ64unO3YaPSwbd8Ak5mnnTR1jz0PrOT
4LEd3AqOae60wNj762pYx3NYYpNwqbHyixp5Q+hYbP0Px3WhKcqN+Sk+TRXECioLGrtr+iEr+f7s
7AlROBj0EHIvzoOGrZxO5kILGSvujF8vNqf2K85B3DuQMhVZok5sv1TIXtsNOAD93h9lm9mMxS05
llZAazJrm0kV4sIg6a1HtPYJF3xQv2ANRMcRJ6uSgWE9RynbEbisGJkz2pXcWcvP4lgH5q3XxhRp
b+nwQBUuiNweJ2k4VJSkdMQVAiSOmcESA04vKBx3gfk9dKwWrfPV35MlV5x6Ln8ErVczZC8rtR0P
cXHCYmnDh5NLZ2tCA7WsQbPMevpG0u+2y3D5/OrazUlMlwz2WpFhHpw3hOK2e+6ehUOjN8u+3TBb
3NGoQW6moRAOcAWeQ6M60D/lhpbyMSKd3f8ZXJuTRbfPDDr5kY44+YZb/TimX8cl6q4HPfgxwmy6
uWrimBBolOGqNgpCZoLPcUGhq8avKRKY6fs+jIjATmValQB/jRBZbnhxLRYZZqRAdvQUd1RDd0jk
a/o0pk0/jjbxKujXZrFMEAflriQNh5j1SwllLRDRi+8wsnf1XEXXSwHyZo1RaGi3EoKvV4vad7yb
K9PKgDkvhi+MPFvYKVuY9h3s8yG7/7Y6FLP6fWy7QBIday4RwTnZxb6yhvot/wtqhlIENXSoxX1D
5N2B+DLUnrLXfQbHoFX4jBh6uNgz7eX3Tyq2lBWVnVgepW7VqIpJgEevAA0ltRmBm84UJv4T/oMc
rCVIOG+75pq1ENfMy+1PMtyC+1Ln0XhelZT5YN2hyt1yI12cIief0Q/HnHJ4j4odYw4AY4iS8odu
e0UnUunGwZI6epEV5Cj/J13rSpF+Sv1Eh+kuyLKKEbKQ0S4Nc9mJcem814Uz3f5tfFeSxzSQ/WbQ
XhbBLD4zlYL7St1kjNAds9Mx7LMqfVj1zX2zjX0CqsJ5dT1MmhdHQI8AlXIQV/LV6gZUdfalPPIE
SDLdRMdzFMNOazd3rkg1mDQm7BcoNOg8hXwxrdI+SIssv/n+fHuPeDYvYLlyOtykDfNPIERcxHuw
mkgL01N/YHpt+h+yY5sRaCagHAPX4sY7X0rLjgVcAWP5QH5gG4d60cqRmA9Nf2aL4yOUsK54xCki
cH7ZT6IMoSU/YYxxfSvlH0N5yMHHDVF24NbON8jSlg9XXvdXw5I7ytqbzjGssGLm2nI+7k6Dc8mM
o/6+n2SQ5ngZljk1Whqaky26z0lU09YHyX/CL3WNkVUNtL5A8u5Q2y/LUwdQ/zFwhVYbyt/JtQ5x
rCDj8EkTfrSMg6XqVysEy8+Y/ddG3+59CO2sleaJXjr0HzCuVI+h56I1mY8/KSO40Sk6zPZnLCR+
X+K/J5DMNpmJGVwAY7FwmXwSeeiBmuU06xIblKdXIojMawCPj2yuLNIjGrQKrv0Kd7YllYOYDkzT
BT2bQhFQcUxQdX6t/ZjPXfcYN7nR22QphjX8oQRPQNpHmamAYaIAvMIzz/ttfUrDcTmhM68/msW7
+3z1eSyTLQRRZ8FcMTGKRGArzXR6GhvQ2eGxo/xz2JRJs5PTZkTAqxZv+Jh6tZO9tvjvs7I8NuE6
V2xjAtP62rc9TvIuIdJJZ+XwWXQPZNEE8vymAB6mhvB8tVDnCnyIe8643WqbO0Su0QMDrqj6rdB/
uyJHJWenmbhVR+pAFJ1HORM63Kis3G3yqQHwXuCN5I2uXqP0GDWPGm2UqpR9W4myylURUQflBGyj
++OofQiQcT4PqCKK2Ritu1tr8W1qpDWktNmp0vhW4/o4N46UaTW6y4R+SJNnX3Du3cTr8cdjxskj
9gvIpBhD+jEytVZGj8lkUpqrB2ylhr0ItwZRxPby80NT9/udCUqmA89eVFqnrJJtrPT/NVFyxRBw
yLibc7wju6CoWCqC12hznTPHc8qk5+QX7aqjhvg3HJE2v7bzybBxJL0HXtaP2JHuC6wQUKAnqIeq
DeK/Lscwj/CQeh1dA+G34YnAckiRdVxNuNRbCpI9JL0RV8eHXim8FVGIF4zCl63SY9C6XHF3qz7F
ge3T8gtQDQHkEZTj+smWoH4zTjXkQR+QAuGdgjB7qedpMu86BTUmVCkPY1WdnpF5vOcaRVG/zbJz
ISGA3cb70gRrPQ0PhLydkSYzY8Xfy5aysqVj8liaEnURY2rxLaATR+tJ2UimPmIA65bLSm+DATEB
zAWh5PyG/JpEzdchr77274yDvMhwPldJ6GMAFHZwAoYJZHdTYGQJ8/YFmPXqHLFQOHPYExZ7aFyw
imdo3GI5pUaKKlbXkctoHAEg4m2tSNtTr2n/J3y105lcJBLtX24H8qey+ThtuTy/K+DYwafgqvWA
FM1aQbWCtCSTiQwPx6C/koJojTZ3ewQ+aw4j+4FRbhmN8K1SKPxRG321Y52c9J3CDRZcXGR62N2G
ppqWnXRP4zzr6yUUstHF+rfj0hz6b28lysCtinsbudUQ16Sq5caMImBPRSano8xzud5ERZn8z/IJ
L4sX5UXEwGt74HFRs13lwyA1QoS6BGcqmJJLQImKWEqAgH8Mk+1YTk2CI1GlGxAbbe/t4LmFioT1
kF+u4JnkToR8+04q0V3v5Qfr2oz/ZXdBBIlN6m3X8O9r99hz1Xx9mIcEPY3ln8Eqlq/kLaI/xBPt
S3spmGuerl2JJshxHbYjOWubQRm4DmOjh0V+X4e1OFg0+Q/FpboA7RHWU5u9kMTDkJ0dqtGc+2It
7w1Rs+SjpO6LCV7HfB5quXY1jiH5G10wlWXdf8KuU4SfZiKKjkEYcm6iYcTGeXjf8QtQorIcMu6r
Z4mWeyLTikMZG/UtNVhBWnJ7e9a6kJsQAYgTti2GzPEstgLPp8wCERgm2gs/ufxnqorxpv7gAFoh
JfLoFyjcT/xgcds+vFvwb9KE7MENEIh5XM4N8TcqLSIcfKj9tpKwSvuFwjWcieK+cwGMV2qpJnVB
ulFrm3ZHeIE2ygIw4jJiD53O5fLyoGPtMNjIOGvUYqooM7l+schXp1Bq3I9qNZztl6YtrvIXCiCl
AlcLwmYcxWRMMT8o/1SIgK1uH+MvjBlN2d6CgC5VBkmD7RPu7JUThB7swjGXvMY6KZ0gm/WeH4/Y
yt9I4EA7EepgXeYF7He/6035VR8+I2c2vWuOsIi2rRUv04HJm7Rh43YJPdltqoLAdlVKVn87cd+2
P1817OCP9lCtpimttDdjGlKvNmTzbIjxEZ9p7ePtOwXNbjbXpTR8yAIjU5PyBD222qyJwwm+xr2V
d7r7E7ONuaBbwcCg+QCWWrCMr8LFII59mzDKHIcSoe+taIUpegxrmolvWVnB0wZzw9/lGiD1KeJU
LNvHYNbmrkRFuS+1DnOUlkW09ZEaUEm2Q4WjF+z7VrXuLp3sy5R2SrHjBsKx7NCW7ICxVBUhBfhw
KIBJHoD2Smj2kkhiz8xQ/2f733QGXJjfS3LqHGG/EFF6E3e1By5r9MPCgUic3KL1a68kRbwuW8Ke
C7dZHxrblLzk0+UxJa0XZpAu/7SafIztxHbmyseampD4qbZkF6V5gBqXEhA74iE2uzcw7F9VmolQ
wSWb5z4cfAMEivDf/ENEuPPjfP111DzbzzjQfKGh4tnKXNLGiV3Y3K9o9uhbjLfb42KBqHVHHiCW
pR0L1DOZdPYm1WZUSwYwk6N0biBc1qi+yPwSbPGbu11TUqwUwdQQ5vNMLIO43+h0maB7ZiVFhClv
MHaZgJVNDjATpgUFDXDv0QRwDcdS2FDxn8CQBddWRPZVulFhy5MPwSPsOxN1qdbybABNbbg3lO2q
6tnjU/4mG+BeO59xJPwDBb3N+9yY43ZIP/bchdCoebqVypKxu9cMfoE33iik6BlMl9lXYbpbgvsA
oKa86JE8YiHjLHLkOtL0IszwciUEc/1A3pDL3Wqp30exHE3nF4fr960tuLkEb0xTxvv7agjWlB9R
WSTE6SURwc8MMXxOS9pcjyGvpSGfl+hjMogjiCEbElFzzbJeo1RFdCH5vICn4/gvIp/c3eQtkFkA
dzJMH/N3b7ZtB8CN7b774/eJbSu9CNW4fp0bpttqeA5wqOB1fO3ozJuZD8EA+68TJKJGMuSpJEja
hdcJqV9TIgltV7L9vUUoeLIRwVt8cy2zq7T7Sc0o1i2xksUBo5j2Bg2xIM/PUoimzAP6NlNULYdE
2TWaj2eTW3la7vOnt5YERlcg6I9sBkxgCMsKQfalhhRjPUHKyfvC19f5I49eIMzxuCqAAPjPrjUt
jBLK5Qq0SVRQklmsPrVPej4jNQqd9uL1r3von+pEyAve95ICh9epmt/afiNK5h9t+MYwfDQHFF1Z
IE9rv5TAZeCCG3jKHm/k805xQhbTkLy2kaNsUzha33Dvv6XYSOT0Lv5kQ8lAYdAa0oGWiTq/adS8
8UeRPnvdZycq1c7TQhyJtmhpvclGoedbZRBKOgI709r/ZHUZ1pstc2Pbme4PrkdOHU492wEYa6pP
p9IyfHS5rhkkXFfo+V8BL3JnbXmGiDc6YDyOImTLjaN2sL5eCwYnbRrx3eq3exoX
`pragma protect end_protected
