// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Gud/YhmqKEWs8Xd1S1bUiYBAb9usH8ScUqdEp4Z4/C8fzsO9YOvkMVg48W00BTl4Wz7G/YC7deh3
nIhFwqzZXPG6MhFuBgvKX05yQpyCnIqjyMO1JIzAvIYNwhlnZzxW3rc8NELBeBxU9fpM0bRNDYdi
cz/3pe3er/TbLqHRuJhxP4gzmL2aShJEDzie15NuydlhNE8iJ/7kRMERw5FNeqr5hQuNJguYWtqF
jgG4mxUBArWqtaFx5z4iHIxVq53XZf7LPesfnesC79OWBXtcL4bVs28tokU8/QK4Cr/xsxoh+AK+
aCOpO2gTXvczKJhfZSTQoTCaExQQohSsnSlx5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
uyyuTnNimaBWqvOAJSzm9p3fBOqf7aa7fCTPEqwtZHOfV+kBXUcZBP8cyE+8kr+pBwwPsfjgNpPS
ebNzcfZxmuW3z8QJnjG5m/KUGnAzxKt9lw9ij7jlU3czK0GE4DBWQ7Bv47e+vq8n38GFpggAWb/n
WUbFX6kNXtTJ/ECvylWx6eV9cOJqctxKGwOOm/kt9yRzxQC6OoOwVhe8ULRQvSTJ+AWDE5+TbpeX
jqg5rGY1A4QdkZZ5VbW4zi/O7zbpgl5prD8qUgZXlI/lZ/u85xOgdGDWNDM3GPU3peTZeIQGVdV2
RZrWu+wY6A9G3B8ojFXIYU/iBF0ODjxs0RLQln8Xh5o2tpu3+VTr3VRR+5gEPBjzAsiptg9/NnCY
7tMh0HGSFYVIuCd4nZnQNuXpXkq5ec/knKDW57y9tAHSKbLkzPik3DKvycDhmhDZv6pzahAP0dqC
wnZ3WkMMdUgulEfBNQGYdMnQGxCpfwTbFIVurS7oBfRYT6kSfDU0GU8B174fUg5+U9Zt/hZl+fTN
m/iddXkpZOGRbKYJVUym4HfUrVGz+RsOMPDcNT4s74Nc29YpaWNRtio/+uavcC/OClTgSPb3ICYP
B5P15ECjFyD9+2ru2QeINQnqpNm6Syb+d/r8DIloJizk4vkWJ6JKuYZbnEzTHpeCsZx+YdSYi5Yb
e6ftBN9/Um+c3Bht9FHJmm8639FAOpz/+X4w1i67X6UhthLYDfu1IZO+NeAlT6rJYExDBHP4BZ1m
fPgpO3PPG8Ce8M+nzK49r0kwTD4Lf5QsNP0HmwOv/OAEI2E88PbGjKXm7Yk0OQn0H07qy0oo2PmE
AK5aBmTeol2PVDFDFIPXsPFJYMp1skjd7m/d0p3vE2TWyrt93VXG1w/KarsUw6yAOgn1fJ3cNeT4
41RipmWBGqQaClAnp+3L83kZPHK6di7niLnCrJyxvuIU3ONLX4V9+uVLDu88vSOn8o+ibxOPLJ0k
ut7cwElv23UyyyVlHDurPsMdHfwhV8LOWzXOU0AlAF5GvmsRCVR9tr9FgLHuiC4lGr6kEQDS1J4i
aA6gj4R0K9HnyxHucw78y29MVAIq3YTdTD2+gYrmTjDdPUDY9Wrn29FQUqIQ6fNTmqFENT0ag+Ge
0FgfaJHQLGCvdMvRU63eQB97xAkcBTfjDmoSqrifGLuD1oa3/zCjGoeWbnegxbEVw9Fm68gDe6CM
x+IYp9gjTiikbDlMCHvpbMkyCrdIgm2wUs2TcCdCyF3+8Fh32g1nYTCRgIeoSZRlzTAtz8Oikk8i
i+LiVIAZPQwnBDpquOQh57l1MisnJJwbi3PzQDybqPBMGihgkyakv6qBtdvUv6gdz7YhxF50q26O
uvkC7Cvn8OeuUdT/ObZfbrPZVIvu8YniBsASsXyQB+Hm08jdrKSXtIBzkqrTASm3ifpCdqOEPEhR
J3M9fc7pC9tsqNkq9RlqsDTsgSiV/kVfRPFRyMhSv3QYTKjhiLIRG/K6baFPBZ9nhsjEY4YFTYkY
EQxTO0D+bOFRyO2aykvDcaAcv0L59clLd7GI4Ve9OKkoF8k8R8om8SYKuUNktaRuiKkBQt7oYr2X
JMl7bI95RY3tpYrLHglXcykpxI5WGdTdySFH8ECEGbamI4sQA6TieGmYG03tHfmKiNvJyeSbCoAl
kP71tiH4bwPkVu9EPRegwAIBLZVE56UX74U8Tub69mBxm/DcqS0UqNkO4eav24tcb461wsBs5Zki
QB+6rShpObUKgwE3c+I1OCHVGckJpLlVHBP1gBm7NtI3Pd6RAOO9qx7e9G43tcYvVnDEawNE9mZe
Tw92OZEGwLOwlpLZYW4e9hpBXEfTGeKH5NRX3iO1IKsKgmpRxGrsTXrBUITLjpv2WdqbENn+XADY
mPwVmfCPsYXQT2KMq50xOvvEeV60eaxJGFtTVzf1hTRa/VpwM+qn04ZtR23qmtpevhDVIRQDrUTr
ol688j/GatH90YtCmwl0do+lZnuozffeRYGUhVehV5D78mm43fdw8d3QDn9mAdvewDLVHEzKmrle
M3DVS4fn8GHJQsT8+g+e/gfTN+DpBPaInSFrLG50BpTtOk9U5S5Sc2eTd+y0K31leV20DIUS8kW1
2PQ6Ve1e/OXEIO8QQTA79tN+vCRwyi3xHLRrv8ETmdhSKzVqwLeOGYCAefHA4GfqRyQoMuId5LRB
qaVsszD5qPWgRWJxC/law1MzTV4RnpS1vwo9SW0aRvlk/dSA+F8zyaDFARAnrEJDFO9LnFo6sTzH
w51yOL4yTphOLDGTW9TWdHoDUKA9nw76YBXe8V0BBuGu/ShVOfRBJhLcYRjk/Kp3ubPrvtBfmFMZ
TDJWVWT8zvFJS2Ic6mV/zvpA9gib4G7SUwFKoXFz58ZUCG9lHCFbVZpCkgjYnpHEkIeZitgOR7D3
13aOlhJ2lOKCRT//kFzf4S8US17Pb2+1eleH0/iDG+kHkzadON/z4/6ToBTeEzR3ZmxHy/qMtPM+
ap5VXAguZBlXI4CHatPVFX8RNwgoputekdbzRzKoOy/nfdqqBsAKE1mhNA6hv8JxW6F5NZi729sD
PANUV4lWeqCQxbgG5ugHXDUsfbGQl1tRzP9wof4UkcGWZeH32AcY6Noy75oXPJ84CCrBK+GVQTZm
oRyMo70f/Wte+xMQ7CIt5+PRUoKtbmvdV5Ny7cpj7QhOFEm5xrJtEROLP21l8Nf/tBX0QNV8aoNh
TFHaJLXACUVXICnhIEjCQA2UGyIVsN6rlmEUjkLPhAX5Pv5Cuq/2pLoJhzLQ9z4gf+VEWa6Euun7
wCErmY7mc8eRsHjGrxdX1kBnwLd6jQZRQ1bRQFmfl981oK0sjC0AwZX/nuxUQQtQjI51yR+ySFTx
dd7afvPWmYucjBHTQNGxcajb3JbSDYffaDZcrnB+DqGxEqlIyD3en9W9V6VSX79WE376YzZMgQ43
BO9LNfSQcXFO7waIW3DnX+hu/Titfb/cI/KyD1BKgE8/FX/1H5d24ftAae6KD/8wm3/hvPolUcyR
oqmHBFUQTfiLXED3RHcsW+NgikK9MKI/u7AZEiRiDfWe9LZJPcPHloGjF//YPeJxUbElUU2ZaRxg
ZD2GjNLM3WlQHjXDa8WSnPpioSmAbb1HWTIYDF1qtKtGWgOTDCU4NDIyN0+Dg9uuEnbMBbJ0CAH/
bYI6xujnVMpIpwznDkBtXwt19b9a1EJ4KlYvL9hVXPbvYTp1epzPqxmUOKW5QT4mZGWKRM9p44l0
qDs7fXT3jdWDH+hSpP8/jYBt2PPO0E2ls9A25HFvcSKpotMW6eYS5vLYzQixQJYdevOoP4utFtSn
jvBz6yoRwn2GFQRa3v+J0Zh4wmYKytbtOCjXXqtyp2aZQu3/tM/YiCtXiebqU3iiGKHRx1L2pQPq
ToebTdFpe9p2FA/gdC08uDUvM8D1scl69wbPUSDKKZPk2JLG1iKc/MYJbt7tMvIp7B+W7g9iKaTZ
j9HZ1A39jFi3B5utx4xROtI4+dntRfwMZZsZiOYKTEOuOFoHV8r/LJNrUuf0i+5qct7t1ojBmrnN
H+myGSGXto0jJihIYtDVfS4dGSZW687jvcqQl8DI76g05rTID6jzmk0Qgcjpp6sMRPhz5Esn25fK
2l1hD7SyrFZtZ4w+mF9Cg1XgHqpx3N/y6ttHeH4w1xLOihcUGsCMr9OpMzgYAyppXP8KQkuN0Moh
d/8UPkoxxklXTmh9ryV1hoPKpiVR9zY2tAGumkBR5A0DD6fA6sjrwWnSOyI6yFk83ukfGxJZhpPS
wfA+QxscRE9Xj//DstwHmjImXFUVPG9WmKrnEe1rEbqN14cDy1pAq+b20j8pr22nvqUzb9foCjL2
GcVEWEgfpkzd8ohVAYKc+FkwyAnuvZUrajTvq84GStOJq6HH3Z1d1NY5MwAv9cx1NxZlm0GZuiIu
yiwNuA97tpLUsScDgLTraTHz69PMggla4is1H+hcHE0S99xiv7V7wQYmJiDXxaRyVSDoHNRuROaQ
gu+KqFwzGe0V5dIGr09HIGksgyVqQUTECUVhEHrtw++0aN/IWuEyLlX8xOXSoOxqRc0sTb5YsosV
+XywIvmreV86OplCTpPs2qXKBacV68f3jaVmPm+fIsRAlPjfsJE8COZAasHx46t3tPThQ7VHzngY
WGYPH3s9Q69/LM4gE2qu/hBO5a/EE2/Mzw+IEQaYfZDX+W25D/RfGNXa3cHzOu0qrRj6pPRd9zQH
bydDcWKsGl8sEOiu5xf+B4JDojtomz4iKBBadHyz7oYkis3iLo/+NTcgBGzHltNerjM/Ow6eMbpN
sMUWn8enMuQ/AcLLv8Luqy1CVUlcM4uThRvlGb2rkw6RZWM/waj/CRsz5I5C+d81E3jR6NS7VStj
iioRQvfy3uj+A1guvZ9N9gwHKJFSylVLgyaMK47Fbtr9wFnxpEYq3tw+BOxVq9jiuTdS/SIbVDO8
ih1/LiB+pJQrW6/t98W78ooxqnoFo4bhx4OiHPRIjLxZrWr6Zw/nM+ZHHHkutj9WDMpqx31BApau
ona6iS3CKf6i+sSDrkrg8f8CTMc92omzyBoCarwu4jaTG+tqnwHXPWU9Lg5yzU9wMlNhWVFS1Gt/
HtvMHDA2g0dHVvXXHbawU23eJaJOdyLjsRe1TBOrH2jLFluB+nwvdWSP5v2jPIPHIEJLNvzIkWxa
/YCl6VhykDIkrtb416z4TfwEATMdoIFwuxJmatWiws7MYYIf2SHxRjbDxSSAr9S8HF2YLhlVOGo9
bRkzLYZC0qQrpltccb6F0VUa4XtYFMBstN6TXW2LZtPTFL3VG5Qm1Bl7S3pCSDVJ8CNzbWYpYYil
2dyKxY0aOmi4Twm+YyXb5ac1H41ewH2Joo6bF1mI7DuJqQmufwbnUBuRp7pCo3DMkhRDjM/zOXtS
kb2nFqc332dgnJNM8sMBPWlXCgpkjK1Hsy2QDCfu2fP/GyxTkz1NGbVrBnqIwJm7yr/SSqJSygNC
doECg0yu3v5PtEMDWYpO7Ct3rmw3rGgwO61OaejCiU5Dpi2osqxQJjZmKxwkgL3HvDY2wFmNqBRw
dTW0ZJBjCHP7Dnp2lOeoHdKGVTNfNBq39rNk++wBNrTnqNQmLGCUnTRcBF37syT6f2VIQs+LgcM4
L2NoA6Wdgiv7XXwiDAdJplHa0toOCQOtmtztPfiOZKXAeN5rbJc3FaOlb35OS48mAw350qOYYTgt
2BL7qEnR1dxXpE2hzFM3VbGB5sX3Oll54Z+HgH3IpcACOG/L8zggPyhIyJRVlq87j7ZcAGHdJk2Y
dx23m6T6FoIFtuXL6sypV9pXAIuszg31Nk+eXeUY7FDhTg/ZMVQomtDXmv5Zn+Ifrnrhxbwxk27c
tWNAfFUuPajwYWgJD2OjLo5i8gVzPlCKdMO0W4t98FrlTXia5imNMT5YUtFSd48NK3cagtSeHa9h
ay3TcEEOG3UfbVlRH4rLaXGqw7iPfyazL4wDAYnkuc0DkeUhxNpTXItsw9tVAVxRnhhtnceYNPi2
VyEQupjUEs+q8APeD6Ya9/Nk1jOyEodj955elJEmHbCpRKHcF7iWnfdrPAOmGchN3/Hw/7iLNpEc
w1hW1Tk8BpIUQFUnLykAcfJSiq48HQZ4ngw54+PK7qdnKn2x7yFrTx/e8su2zxaVnpo8bBav2Fja
0dPbHGByb9ovCNG64eogD71b91muneYUL/0WqO0HbEIMfidkoe+WJPoSrLP4Rx5kvtO8LnXFbbl5
tS49Bm639CpKkY7YOowDbJy4MXGOAgx8gEnT6ta/Tl+v6tZ3iTpl+nNs39p/WTgiHAFyx8w+rw+v
pG6hBWqreMBMTw8dfN/y61Hmr65GL5mDsNYQQkQ/WETwljEMA8RTLXOEaz7K8Kmp5//NHWTShI2X
xxL0oUwFU7cDhASiU3Aettq/JrfFIo6Mg+HY9EIg+5yvlqGW1950YsV81bErGbNofvhGfixoD90O
T4iyQmxhmFHmuAeMWC8vh5os7ZqVH/PJZ8vd0g2Pp0nRpCPFwGZQ73SPSpUdtpL0uWDVki/SDz5L
6h7Jy0KSnoi8TQ/vKzyRXOmDig9oJxtnxwjrI5s6G6CIb5lvxxvqg32euz1L6kcqqheT+dKKteU4
WltwaOSC7AhGICpHDkFogZhI0YOtTX/H2hx5MM3VhVgcru2tF2gZzw95l+KfbmSBWcB6a/PH/snG
AJHDnQ16orEgxWa1faGpXrD4Z8oZeYiwoNc4o39h65U/EIABP9pwUskxjS7Jy6LWE0K4OuJShrUP
g24D84QAgiJIxO4tS3YGHAh9FbIsX23y70P9+fRplL7KYxLrYXLvfeNrCJnUphGmHfNBWnJrYmvS
4TAb4OJ9joIXpLAXdFzQ4/MStcENCD6VFek6c8m9carDt9d9bUE3j+B9zG+Sncfqh3XrLi1TVlab
ap5dfR5ruQ0oRUFA+/htTXE4Tsga6L0tcirx++3I5CeZ2LiqcMP1cdWRc6aPSky0C52foF8qiikX
TQVkcYSTHCoVo5Cv/xCwOOHfAxWTx/z2LRFHRMAERZWE1+fXkxiYOIL1vImLGldn1jYnq4zlPGt0
9mgt9AErjRBGBp+hhPS8VBvQQrlAgKacQGxVOpOjKvm7NvJeoDjAqFvz2nJAdFtwHJHZLBrXKg+f
rgzyeGq/xa5RvfhutcmUFEKMBF5ir41BHZcqr4HbTzpcunsloYsLBul0B+UU/V+/FpO916Fecz1j
rwangi7xbB6YXqPQZbc7HwmQSwrctPL+bc34OxSoOno0jm6n993WpAfSp3G7qZJrnBFeHEs/Exj3
0WmwYpYRfAwaQ6Qci0VifIAFFkWGuWQWV9l+h595CNBlPjfgH617T0H8rCpYnQHYx0Di20XMjdwt
Vqv65nDwrxpperoqlEnimWtBh+q4/NcFjC1IrMdztDvg8cCEBSplkBvfw/zRuFVXFUrshGfcpSZt
jew+yfMmFZFuKIWU5ErSjkZGRxOmfAftxf5XF0aVwN/8KMQ+3sNwAWVMtM9PDLwvZpCAvOzs8lTj
R4StaGl39+YYBz+OZXFCszZG4JKedqMq7Ad1hKMAuYDGlNIW+4dLSEgCUox6WqclbobqXMgpknhd
7RixKukMAKl1E4orKO0NEmaXsNzXD34UiuXRq8r3GbWv5g1T7dpS3qi5p48SIeQGVbHiaQOgRgcE
LEw/facBzLD48EXxxmcm+SnnZ2at5Y9TpY+WsCPEltGF8DHAR1Z4Bmnle4Ev4dM0BWMLIamvSDmu
6cUvgVgs3Hsv9BlemoS0OBNa6m2udtttSDLGCG0oj+Nj5LYvedHMWdmpQNKdWzjPimFKCT+gtQt4
kuwgTwg2t7ejFaDVplBuNb+7LZLL0HXXyIOU39X3TDuReXwePZzGtxaZXAhUnNcZ8S9YDl3IrsuL
HLqWrocAPcYTE9xETNFiOyHuAjx//yFcu4QuLlm03kpqO9kn9aTPRXPc/cD6Dv3F8uxdXLlAqwt3
HFGJF316bzdUxB0BYwa2Zk/UmayoewOtg0C4OdKCtr+Zc/Xir1AFxMl0CtPmRZ53zJXDrHzoRxp9
IpbX+rKKaR+JTKGW5KdHxf5XjIL3kp5XaJ7Y4ns1OLUy3Y1Qe2ZAJaaW8VbqLAFb6rrBnauxA1tM
v/ntHUXVhEjbwGzXdBxR3Yqlu/wlw/QIwGQf1CDkwLxoJzp6r6aarapNhwyBUiuaoNuEDryikeL9
5CEnaLBGHm8rMLXZjG6JCAaGIg6mL7zYVIH1nnHtLvBc2SURh6Wz1L3Hus8syeqyYAQm0Q+ZIcka
Jg0uTZa8ps2S0rtMx63eO0DyfXl4FSZ35ezLY73uw1JngvNIcQ7Y2YoQq+XiLaoL8T08H3o2nl5A
e98+g3l9TlO7eMflHbz8UEiMLY9yJ7PIp9yyZ6kfhA3KTzXk7oeUssYCwoO2F8aYuXqaYdlwl8ld
ZNaQRnjpxFlcReKsfH5SNB3UiZybNgknPkDut8JcdbYlxHv3HydwVrw5f1SvitTt2xsdGdX1ZsdY
JSm8yhpX0WDUvhl4PJVRRHG7tQOA4qNFAQQic3DpAYfV4X//RkjAAkdOj50kT0O9FTNwRPJyLLI4
j3Hs6HTsuhimZs3wfXLEpOLqJhBU68ujaxFXbscbOwtgwqWC93u4xunjdhpk3iF7juR/d6Bk7CFG
4VK+trfvRqS002q1/9v8vIZapj5qmpTXDcWYcnuvWoZkiYayqWoFiXUHT8BnHUZR1rfEoion9ydW
WWkRvW++ZLsriNSUTyVA1vIC4L2eWk/2dqsasel+F7ZbcV+Yu2rSlsciJoSdGz52Zj0GgHafRMiG
53mthTUn7WwKtUkP+5hGqwCf/jBxCTz/hJNlDRvmBeCI7HbnhkpXRChwVKT45wW8M5h5rHY7derE
Jgz+hudbOY9FIclWNUd8Vl760hObHU52RsF213qN0pKzf8BXtXec0ALYI0Kn5Z35j/wMW3wGlFsZ
jxFJsuD4EXsLzs1UixJcuf1skIDmmbA23mb5H5RoTLk9mW4SxcI+UvFVMRkkInJRHRvfBZQqBNhS
MFl4zRUq1xX+arMGqWO1IiiGO4inv//0av80IRLGWnUh4SoqnzNWnbWNTWUjPoySof1TnXCxvPds
p0mlSgvwd9dx2tShtB/BzlRgljMA4ayqZAMIBKKMR+Bmr1+akULv9YYIiCE/1dz948+tMRc9UJ3g
heXrfWVsG3SVfFFzbfgyMkPrDlBIka0asgRnugtVW6iM8XsScG84jqiT/Te2msVMjM9UJIOK1wWk
s4vUMppMjo2gj/HSY2zn/TxIaXV4FkcpSnc+Hzk3ewuW6tUp+8eJQ227aNIQG8cpF7JRCQJ3pK5+
iAhiQuUrZ4Avl5iyf0VfMFKfdgGHQh0STFNORjeqtWkjatLeBmpzF9+qkbFRMqXgN+uUKasnxHlr
7bgLnBpKtQENzaF55jDKZPWS6w9p0zrdYEL8Vp+i6FQ8xKwIxwkpFGfwyczoAkxIBGnk4AUM6otM
znxFArIRbwPxKAg1qyr68/BBskk6yEyeqWheErmfcxpwLhu4QxSgwqFllNR8AQDSvmuq/2YYP1xT
QxmA5BFjnVL1VSvd5Ajn+ilN4WzDWPVf+Y3MCrVWsf0rMJiaKxq9dcjCyqrPHQ9akIOhy5zORKrc
b6t8v1N4XWJhsjY0qh9x2osbLV1bzOn3FIEmytAZ/QgM4M9pvIQIwD1y2Mph0z19GnvEsp1mpkp6
NA2WSzGB0KcOp/w4QvkF4jzFUXbWrQCvblPuADypgx5CW23o/IWmFBUvsZsuxI45bB6aUS9ezwFZ
ODA+zLWdmCbvrz3FXMa93Uw11BPauN+2B7EZuOc29GFOzshPWAm96si9vE6wueTgF8FF91ZFXWTt
4JTkkdcc7O6r9tYiBh3+nV7oaxI8lDhHzEmEKOdWdxXtZ54NO1WsHqM8p61GZGUZk46k7fhbvsps
cGAN9hWOSchmsHnc/xywq3tZzad0inO+p7bN3/kH+BOUAIpR5ntmDcbWSnGJd07POsbdjvKmExj9
Wg7/A+GjyTTrblW0LaYRnx2GCAwMG1nrDyGxdrWGUDSVp+HNfsr3n0tDjDd800+5RAuH8p3P++Ki
HhUsQJyJ1ZCe4/k8Yef+vUi++3S7o7kopgsjwIdKzrO7FoQbKZYueMD84KJj48bJ6OJxMiL8PLJQ
ZKPIcr9YS7YmuzMZC/AsPx1TyD06ZEkDvRuVxmuH//Fa2VQatMpxXtxd6g51EfpDoAxEgKPwPTsS
i4Re1YcvGeltVFwiMJFOT4DvCeLjVPzebkEvdzI9Jbcv6+BKJRiWHozi7bbYJXbv/sYnkzmW5rOZ
aKgysGzV4WXLYdyT3mc7rEisS8pl0xAH+3x0rdFkgbJJJeXQsOwZv7m7MSskrPmu2XNuLiqdQYn9
7KJgam2o2VJUH1tW/MELZcweNzU9sXHXxmd1bYfMluWimL74HaCF6YqveMsjai/MN38eqJ1NTIVX
PeZX+JG402Yk1uW6Gu786L3JybZZL9gTdzyAzcSFu1Qfh8dyXJS7ZpuYKDCXq5qyybN5uMNDin38
bR5wUre5mkTvMj76U7C5W0l/N68Yx7x3HoxqkVFN1GmGjpB7REr+AO+9RZmbtH5pOHyjvjRN1GFb
C46y93UZ6ooQs3ysmZtOj0p54KW/kxKrDYbCYtEHY1xEC1iG1Wue3EnZ+jslHvuvXcWiUEIsFvjq
OIGl7zZSR1Bn0rx1m3uX9KntPoeNGf43fXa4EnQ8pG7EsOMjI4xxEs/ZNZqxoKNgzJxbN/gc+pVE
YHsj8BKc0xmrhAfgEgtpdwEfD+jfwkHXw06LQTCK5S+jA3A98lvXwozsyLyI/koHOFvaHVCXRSdy
YUI1sA1mLCRyYTsW+Pb6KLcjvaX5yiCeTVsE4pzHOFSEczMHjm4JrDDZw7ajaj0zBBUEm9uIWrey
5EczoB0rnnsPHiRr6SWe9dkkRuC2cYpTH4kbzOWsb1xKYGk7VDRW7xjoXXAdlHTDh28Q7TpjJwpT
ePfov6+uJG3l9QdFI/R96XkKZQXR/LO97oP74F41bd8wLSsbeTUM2azyKD/NBo8rqSLxA0GAFjXS
Mstrk5iQhI/FvrTSkVFRoTJfiXoktQu/FDbSDSDCikRm2D4hmYcqgKNqYyq9ouWGxILDGcCIj2Go
9/Hz78GUhfgg7KsIj5vUaZP/IUdz0m2c9DfEbBpjU8E4kMvfFOnIIxhk7SYh4FUsrYerzjcKYtig
j/0kznTHS2/zMnyFTIysvjINuZghQ0mS0V0DC9NJiOLxuidiheCKZ4vt1WDEWmPQQ7HLZWU56hAc
TLB7tyYvzWwJar0xjzexQyF4Q8GrlQvVW26iPp3v0qTYzQK6ATjSN2+aphrSVV4Qo5wbydwDyUO3
aHropm6aSPTy0S1a2EsfgQwqBzlHkF7RzkAuY5NhmEclnDRvZQu36tSApM5s98h86W9az9iQlGCO
5kpG20e5YNde/fUQAJR9O4Bn38KAKGXc5fzyiX3psoJZeUsF7Is2xicLoB0Yn3b5W4VCHd5S3fhw
Us4GMPhaVTtvCB8ExbEfDtecJcPguRcsU17NqTMsJJgCOObu3SDJUBbzqrTBVRqfNX56YuduERW9
AH14eyHg3+/PLdQ5pZd3yyALKnylM5UbiERWZCRnqzesJm4FiC69i8Oo0wUfhPuTPhHshSGXy8CP
00p7DWCe1VskgwnP77t3CLsL/KhLbt6E2RHT5Jo/KlTrGNYCzVk6kb1sc2g8ZA4NklZ7FZ2f61nu
gypZTiOls6NNcw7o9WrixQZBMcegyeQP5v64kAzHBHgz6sS8tmpi8/n61jJ9s9d4jGpWrg0FhwL0
/Pic0EDQrRBy3DtbSz6xvGNBpBkLsaZ9IdMRsHTtbPC467fSgYyoZOALPOjICHMT3tYR7ke7Z8zV
QV8WHTtO08S0y05ul+vJdzLZUxNFfWt9eXdLiJ8Iz+7zKFhNKbsHKdmDlvC+JBaFPGe1CCYx6rwq
d+WWyYS5D6ETc5E67YM9GNPvGJcKBDRo5vwTXum2YFIS8UWo76LCHmrmCfGHtvv2p9LlC+xvlRfz
NK6TqLnx8k/Hhl+eVhUkh2po8sOKqjxYyHo6OyaFsMPHXUIQ3Bn2ZQQuh9FykbSWFEmB/LvFjFfH
MFj00S8nsZC0Wo+JNONqpiMUYgxSvRvFv7Vlz7JfY60IZC3BPgcIhxQUQ+RwsZwWhEltrLqVEKmT
8ZZKB61ASwLhCvRV6+gU+FN4hHiDBjUJs07jmBWqUB7lMXBHQT8YgWz/6YKfe1JJ9XFaTZVE5p26
8PwEZHM0HDwAYE1PDHeuhkbTr1+GLBY4Ps8wlGxcPYfmyCw4pY5CohLgf6bCnM0n/hyVDPPoqZgi
mT07jqmVOCA7Ds0pSbEBCpD9Oq9cW3eMH3sfXFiqfv2E3YnREDxGdzi/BFUvRWMmCXLtsBJti4Ni
cXXws3Pt6ZsunlwGs+MNxTIKFgCQqSnYV2eWvvNuUWQ3wjBGDFUl+leP/f5AvTmmfQLMKf9OvnAe
+ja/Z6OyNAICVPeXnCsavZGEYYSKT1HeSTpDu1zqu4I29Gzj+sjHta5aOqjUEB6vvrOKM+AmOUkb
rUXeGMPF0fI9U88M0JsO5bfdIhFIsTMTwHCtRnNDZAzLWfDbmbBejP0p3EV7rDJlWahIe1ouipTX
SsfGbIMN+Koh03dm4VxHTAOfQCRPlQAR0MyToFEHhf6cbppTfcaJ/ak2ektOBYiC6Seb1N7HLBOK
brFZDPeReI3oTYfu7YVER+GEk4YXF4qIP8Qdkk2oYOC2PIVNB2lVlATlh7hZwJe0r+lbvTmyYVMo
T1djsr0e/MCsULoFG8FRHur+8lEPDiLMufgzgYQsv7mRe2FkQw4cMwOIGjxqkriQdqhGICbq5Piw
6YfpgnsPpjJVqJhY50WN+AFn0ujZRq439Tx/Zum+SrCRQozE6y25IrjwirDE1D/e9enZK7axiN2T
80Jj5bPn2QEnAX2Hl6ZEFFe0gO2LbIiFm3l0pRR5mVemZ3XPr+d5LkCCZnA0vFU7zpNXVuXpQg6V
pDhqd75xcINb8759YbLTrbQmgs+o4TKMzx8RsESJcRpBQcIgK1YNzbsQYbb1N3CLVJptGyKZEwrB
s01z63pMOwGRbkL3fC0BumibaBH56+byOYs4ulRbpFYxGl85Zt8vMlPMoHVw74jUjjNGpejfLzmF
PYkvMYn2vsedBe8+yN3osLu2mSNBa9fr2IiwsH2Y2xW356YKjVEwxjVTgZFpy2HWbGUA6TbKJvde
JM6QdXMx7SbEQPfukvxctqxDgjyLF4JNiqkZfvKvBqwivkkUs5UZMuDca2nj7wiBkarEsPvxUmCP
6zOGxntj3O9/dxvUEzjhHvSA+lt79aIi6ZgH83osxZwoIBK1ZOPuxsEFd3t5lqlkKr8wXShQPZRf
yvEdMy1xEQCKsM6FOrDYsrToffVR16+v+sIiXS5wUsnpYqn+Od5PHDyuEWp+Li8oy6B5YG+iIC+8
py/e1cPVzwQ510w0WsyJMBQk4L6RUuPMmCLxhrDDWuPQTTkYe5p37ozqYF2oMC40NPssyZvK4HLw
Uhl2fs6EYUUwyyB53mVdmD5AqQKffzKx0bS4///btqJ4OnTCQZR5nqcy3CeJFxcu1RPBK0bo5F6I
Iuw6KqR5bD2yNLM9Py1Gggj9X8tWLqJbGJCpam4hldogN5VEjsd/ecXmbaeZXiz63MkR+KJHFSuk
ISRiWROKu1Q/zF67r32i0Yh1uWomRlkD75vsOxo0JQpoGkBE7+8mUv6FKI9UK1tQWcnMVmcdOPQH
zqdbMwB81z0A+/SE8HXUeOhosua4Zu7JGvAK4XigjoB8sAe//cRTiqKPdhqTQYgCFZIKC/AeQ8kz
JoES6+9nTLsT2rMXkXJ/HjFtISIFhTCpTCbBE3fJ5A8J0p0Col55QBKCsJTkmaarYyR2qcM5sc3j
eaqtWO06Hw0v/Z4x9nnHFQVnL2BK9ZTv922xHxxH8N5dj7cBCRv+O+b2fgtKvwjPX3UTbMjCMLy/
vGTvEtXfbJO57mvRMnM4XKOYi7lttbHPhsNEbsp5fWnn5rgC8F7gDWUWmPqQmbOZMnjNzWWo0RZ5
uJQtemHS58qSDe0VIViruR1CRF9wXaAv9oguYIn0Mxm+N8h9i4e2s7Eh/uksAXug68J4NPkLC867
GhRWnt+gK7wPghU+UdlDe0oU4OOvrZ5fPBsbXzPPfdq0a1Wifhi3JPBetoXFq/biyxBw/CeA0Dd2
v4z1qxcUjP7qCCPEKfOmCvf9k65ojS/44k25oDwU7k+r58MjWqSG089e2uGp7KhDmmObzNzm4M6o
BdXfpoxqYib4Ok6WRY8IFW0K7Qo+RLmkVxNbEct0ql1huRSHdIQQdJT/hnX2hpybfbzvqYeeMUgG
5wujp9X1TbVqRKHltfqyH0t9w6iSbQqzywJGljW/HJliQujsCufxRPi7RYsR1Ud6NH/qTfANd8mx
NMY5kZJRFKUx66Dq9IsZHFuTp/NtbDLhYP5OL5EiELhPh1I+Roz1AOT0ZReBiEBae+gkEzJTda0u
7rjgP0p/UjX5eIaxO7RM/ftFi+p+Dyxr9PahDnVfy853uOA7X6+bdLeDXmJ1cNaqBAtJ58UGwIOD
12GYTU01gcpLrdzwBUSI0Bu5/RZgbsdYZ6bax8hvJzL7hDaK4vXVoilkq/pPqdrI196XUKFLp4LA
bwAy2+QJe2lh3eDa+oWKJwsIiUht8ngGommAdnodqS81TPEo9tRq6ixwHUjODZqKjBmWMFMlJiq9
FRD2VbsX0I2lAY4HlBN2tGkyP0aUp6hyfyg4rqTUaVlGGYRjs8HZK9o3TZEcKggIjjR286ZCWu88
jXDluHjbAgbzymLt7x/lQO4E61EIWn/L9jvKtk8VFrg5hm9s4ragovZWBKqnpPjuowvcXBr1Rgis
BCi+Hct8kTH1i/r07ElOpJICqL2MRBoiakDvRfwH4yS6Mgv3YtGYWlhjEVOj6r+ohGzUSVV2V0ha
kOCW8x11d06BuBpeL99RXI86pXXWjlQocwHTbR4UWZzQs9cSgwMRThTQi0EwTRSgOJ8x9L/RNdyO
tX76AwdE9HJ514sqlKbLsO/oNTlyw5QlQl4xF0eFYYJqWPJ1XJvMn0KTC3lGRG16dTKd1CfPMXh1
b00dl9SdtW/JpHgsl/EoKB3DwdkxEFe7iU80yDpcWKjhfMtugOS3RD0fIDnOglbDiIorSjR7Id7X
px1fPnNHVld1yo3Q0xi8fuczpvxbLUl+u70Q2XNA3Zw1pNDq6ogtAjVylzWXVthclufQX/bGi7p5
CAHUPiZpOYQRnV50ulwJ8J9W1GfbYPiA6Jyu0AAckkVomFgNOpF49jrqU8lTBwcCpe7m7SE7zHU7
9jyEDOMFpwKe4sT4Je4hA4lUIWq8pnQF49Iy9ogqW0gkFOkeZ/kkpxRXd4HZnYvLqIVWjxvtLJXq
cbMllTD+TeRaqgEF7Zw8uI5wVWKPBiWp1LmfFjQit6YRZH51Tue9rbanNuDpPx+/RxEzNLRO1Spe
V4PjOFLOfzVcwP0XqdaUhlSnEDD6xWoSL5OYj7pO3Cl0Xu3ne6WYGaSJFxmZEsjLuMzbEMuWt2VB
+5+qURv+TN7z8us7y/kqYh489TUsgKDAXn1sdZPtrW5BD6bUtquG3Hm9NPgCpF440pB/84WCu4tK
ejf/irUf2Ih4TLHWhfZehcZOWmQBReYt8Dro5fnEqhJAtg9+1FH+A/M/zYiviWHXBrBo91CxGv55
CV7DLcHzpVGg9XKbZFe+3TcVRd0LEVElGqlGYAULKFSGqUsm8hT8L2ypp9uhfQm7KKbX1IPfHOva
0tXKPmJeYKVX7w/Hy6P/jkQDOzQmQ/u9lMIR3CR1iJVdQLDXzXMe1Ed+zY3g1MGLgcnicbMmNuTo
SZICnSY+kyOaZnpIrjV2AJIhkSHWpeArT64uat1OZa3pGwt18uUC46oI9pjZRRTAGvenc6rVGW/l
XbTVac/3l4d0GBgvO1ZrjUp2QHwTL6SuPENTVuRQcd9oeiiRPYqblx4hk4bRVVP1gzONnrYr1tSz
CtrHvaVgVbA+H5ndB8wF5VHeDlCjZ0mv+zF1icRvLPDz3FlaDXaq5vHnrKESaIZi0wxKfxrlLWnu
rDPRAxqxkK7VgEsIuTc2RtEQ/Wrg3HrQMlZYMIdeelWI1z52qwRIW0SLnJwg6rapKx8uWQG9xg/+
QRJzLYOdgyVBxmAxIl/RxXRQ8cCYla1tjg5aSgPPmN3ODZnOgW5edQHjyam5SMyGFa1P8F+bMVwY
PuezyKzm739nIkf8D+V41HDcgREHuQJPd6IgipIP4WIhBh7MXy/JeDSuCnyPcvvJkaL00xtoZchP
44dl4vqI5CERKCWcYhJzXIi5J15hrzk/pA6RnT+TLtpu+21KKXnUuzimqXJQFwweIsFfjUghL8xZ
Mt56PhEDioGXPUf/7bchBSIDSSj0lKlpS3c2AWoMdOr5rihPaNLNC5tR5l6dKEPqxGggEmYXVa38
jC0QyWRL7mKd57gOK7B6lSOqLLUfA0tnJNrZK2ehT2hy8vbaOMVfwi/+LbNTYPZR3j9QYTA4m8rV
K7iWx2cLAQ78GoMU46v93P/RLFtrMfEl2RrRpRMrC3d/WvUozZlJimdOJjiUruuzOyzeEZ3nv1vk
k8n9Ha/PvFXZY4sOWluUSsLShGAwQyetZs/zZ7pXpt7dXl125dNstsUCn+eJlxBOgDqSmtBLaAx7
kw6a29ZmJDpdIM4hAbJyluO1otd/3KxYdrW8eWr1d1rMczgUSONtu9H5JCfLTnZ6DOAglal4bWVJ
UGX1QVYzkbqDDyCAvOGYDLpI+d/CYlbgpMzRtIRV+gJWyTazOkY/Ofy3uHN/1cCMlhlFYzNcui5b
drLeX9fPjL1e2JWTuhDiWRDmkGsDUxD8pNu8obwb8wfW44qGMVLWm1ZVDM1fKRovm8pnOp+D+bFe
zGiGdAIFU+m+8lSfJ9RnUBwkJ90j6ncjY5KVHD0mDnLOPrOuVFVvEJ0fPyNGSzy66q5Va13fIgXj
/HO0LzXTg9PTwHfkILPedbYayWQIEMLrKQq8iH+IVz/1S/Vl2j8j9722/Hj/OKYrqZAKAD2ywQUp
yyDaK5/DMID67RHtRXaC8khSDszVcfMDGelXZWESAd4IWg8MutzbYs/dbSJYobqhoQfMASGbAYu8
0nddzEufDstaOd9c0nwFwK+BUocyL3TUcxczS83J+KwNJIhcUvxGZS7VyiZ1CrlThWU1cLAkZdEJ
9oaborp6a2hSN19SVR5YjRI9xDVMmDz6NqLEkNP/OiSmechOWbFQ6E0dTt05NkcgQk8iy9Kv+J0B
uFmv2FqzOfwp6wk6Iot5LAYCDk8wPQ0Tt/2wj5b/suehknIeISmBvL81Yfy1Ui6RQmE28dzyuXtC
wkd/qI6AsF3Rn+4M30QKJhufmK1BujTgg2mkX+vZWSkTrI+jBsxT82HvMOPDwsxJrofsFkDEG511
uSuZTIbVFVYvuao2hL7yz4163Y8NbmX0YmA1UQsjtW+KdVikvkBEi1uvv+EnyAhVRKB3f9Rm5s1L
jLy1Qu1Xa5NEj1pl15aj8clzHGAKlbOKxZSB11zVckTlf73tTK8pIbj48E5DB9IeBKYsPBo2a1Yp
TPLitx5ErrhEqdPnUljXePGYtR74O9ixhgZDmyItktBeqNwuUQ==
`pragma protect end_protected
