// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ym8HiSoNFfzXrjHzdvkYpHh7zWfvQx799NO4xUj0+Zh6rNLZGfb0WkjtC2M6PPW4
8vfL/vGtj514ZODPUaKEsp6zUPrWqdP47lgqkyZ3vpisRbV9hV9shtD37ncoUkMx
nGYOzhoYZJyDx4j3lBxTn65WCF+8KklgxfoOkCqHUfw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21456)
+crHeTizFZaFVwFdKE0U9nWDCijoTFiug/HYajPPZ14PLhGv8+WjO6PW9QKEAIKD
DBDvaMa0XgTO/dfr//6sIQFtwZTjSipk5ksySE4elk1CewMNluEyKFCZWLW3d5Eo
B2ii7nQlbYJ/8UIUS3rzY3Cl3Nt3sGzNPdcvj0OufAH7n/obTmZOJbrIbD9k4rcp
C6A+zigOhM5u4sGhew/n3xmvinwFV6IzSX6wxwly4SToKezZrI2dyB2WXXQoac/7
lrRqs0C0XoLeJodUDK7BLSg1evZD4j1a/LB/XWsfK21lhkLCcFaIcgDnAY4rlzd2
shX0pxeUorEqnwwuvIbMTN+0QSrdSwGkmXbvlGLosN8Vt9o7Y1jhvJxtTL+HKDB7
KYiTQ6nyD1FYWG4R14Yz8oQC++0ysDWW+SQghnPFC1cG5BBAoOlGbVsaAXMwmiYK
iP8ctpDWA5Q20SSUEc4RaSE5hh8mBTnVCmf14z9lM4gBqmzdgpOx24a7uC3XQL2K
VFKPFJsXwbXrWn72SwovZnSvlUwPxsMgpee3a4eUoTkYuCTEMl89NLm14M/hmlc4
V5s8IDdcI3bWUoEG1R9CgnlHx0534FgEDwPCAuR82uE0sDi93eZsd/S03s5kok4V
YPQ/1l0qkknmGYMOvxCSck7OwdTVFYL1EeC1MIZDUWc4CvjgLCZLOLgw+1LFZErC
nHUog/LXDjwu6ZBjdzm3shg3ohTRiNvA5Ji89m6lfgF57gchF5QhNyRkOoVLDvD/
0wJWa/gS0yADapwtGRlZ4HV5S87x9blT163tdIk4fAnn7goIFpjZfbLdTBIspAG7
tvzS4NOn4u2fH+IhDO4C4QxVyoPKu7wWVmIVWgckxigH++RGNkV1m1qfZedBI7GQ
fHZXN6m+AXkuN8n5zXVvIag/l3emh9TuhXmJj/ypRRago1qNGlMX9rnTvzEiXEzc
K4KUqPF53IHnXQtkmFtpVkuP1J93Emf7/Nr/XGbOYyYiyxyXtlJbNazx5F0ta1vd
IXY1YjooWlUCAcGOxueFT50C6xHq5H1GASwBnI4xV/a+aXzZxTcN+wm7FAOal3NC
lIdMzWPQ3vhNI99gDe9DFip2fOCsi3xQ3T59TVR2QUIaMyFOaKK0fQWLp0t7XClS
YrD2usOFg14t2B5LsAgM2H/ylynLrsYexTihrOM54RSj5LffHTZ6l3JUsyVQqe26
PglcPD9uLUUz4a+m6SepfRImEhHNVG8C9tPE9L/7ywu8y/xVRHsZL/NeDD+aMXkR
LCBUztJl7HCPLyQ6prYgGNN2aJ+VmpfmA8/hyR3gVBoL1Ws+BnE8a5GoIYYXC73m
j9EHtROBMKfQQHVOMF0F5ZNFhKYo72ZqTFytWzhr2I3n4ekcktz+2JNWgz1XU3mz
alWyJJ3AoLlAWnvVWnd0TgDO3/ZgWVnlT0RkDRGNV7vAZibiuMRg7sCeXJpltewr
OxwL5vnx/+uQYlbbhhzTtn4P+elZJlQOKFyZZg7qmoBbTEsaub70ZEcZNzqZjnaQ
IjVn7xaROESiURW5m/3f0S/3gDLF7qCQfSJfVmXzS6MnhVFCwGe5j+JsG4Iyw+1J
g0b2efLfj4RKqA5Zk6i3LzO3qT4E1y7rLFNL52ScG5TO9+5Kl1BZKrujq8b3Euw4
+I2eY1BVjxJ52Aj9MljTbSHePx3J9BczHSYkV9+HLhx25zEc4cMMgwocD4HSYxiT
6RKvtMTmIoImq9Jf+r0WbVoDD2obYNkVUE9PCEKgG52JV6JU4pp2fAdAWGp5QXqc
oXTn6cDE4T2E0m4HymmzajIcK2M9A0p0MkFzT7xDUSldLlZJRrGwhMRRbW/qrlmJ
I5aQLeOxvyTtPg1PvRyyviJL+WgtMksUEoydb3i0xHZ6P5HvZ7G30oxN8/oKqxh5
2fp2SRd9q7kYeAWtAsroTXOUff5KDgf82VVKfedveU+zKQCMCwGo+sG5erGl/Cqh
1m3yeF9ijpFTp0zYorocGNqF6+0dw37hEQm6FVpjYl28j1Mh0hnvFTLEKicfTmK5
FpmQWlJQvraQsXtDUBwnB3wEmgX/nat5EXvPU0a4BciWCJz/XN4OPsU5IaY8CPKo
izuhcpIBrF0LQxxAAn5PikzRhX/vFruwEvS3hugJHnVZJb/Ij0pnPDDlA4pfLjUu
NIyhTQDUBqhDTlVHuTQTqkhiw8YgQkW3XJyIe9OtlX5f9dNJlo4aKh9i4uKpCBuu
IDH0cCeWdwopYS1QyUG5Ft+ETxZ61py3cHAC6WDTXdgrx63y7Y5MoEdFzpfUUL56
fciEFLS8CgRjJYyokAEynH245xrJFIU9G1oy3OU9Pd6z2u5Hnnce0t4+nhob1c4e
SHUuB6cobzgylLGKlIzBfuiRFGN4VL5wEVdPbF/8lL+7PdTCCpvJirxfnvf6XZhZ
OMvRCs0hCGg7oVZlgaQzLOD4BC60oiqAqA/7qZa6jzYU8l/upI/sDXA3yTYhkVmz
8SDspFUi9HM81rz7S05elJOSEF/5MyxyhEK9FsXDkbF6VSdh6F2M4dvia2cuuZWS
lq1Yeu5dnDOXouZrzFk8uItDzF/XLsGSw+NsCCXqCjougHcO4ie6MBQAPH07J7V1
PmFFbQ9iO7xwEt7B3rhM6Z8fS2N2S9PnFtsM2rLqizGSm+6joDfPXCoqgKlMCd3o
WSuB8U+m6MfR3uO425mMGylxtcjIJ4NdYYdycFfYdwnfDgUC2NcGHcL0t+z4ZQLK
X5ijIG7N8Crvp437NmZvfq2RDSzUfoMrdqAM0fdwn7Bf2Ts9rERf9ejrrrmVMDUM
CWjx56I2VD8PhttUmGRUWjeVvs/+UCv2XTWGlDslNL4p1EGDvRFeIx7GhkZXODuY
N8uemIwqcVcUmxDbnco73+WB8l07o1ZpOiGKyOk2Z/9me0VBTq+tkSPQf0ATh4pp
eCTPhZMCpBhnkUHwx+RZ5toM8etsG0OZIOgIpQ44LJpVWobnu2VOfhtbOsvmImwk
Wd+6w67P8ypP00M181UOz5QESSHyGdj0pkdCdvYU7+ovxhl8zmCsEEtU6wWuYGnW
Uubh6IyGVUv0ogjY0CVnhAKEUwlurgAGioubUQm/gzlcrq4uUuL+wh5Q2ROqsRPf
9pZ2ejlITJpzkVQh6EBSg9lk5Z9xX7jNtNKU2cGIQwQ7gfD9l5Yg90Bn0BRxKTRl
pM6HvpaEK89tDu4M4P67L8S3O+gqrzhNY9IJL0BF6zDGNVU60dQP5qHUtrPc2pL+
v0wwAsLGBlJ7M3U45lYVLj1O7Y5J8r0VgZKD0b1H8+Z1VogtaW8l+H0kCf4YSTU/
RU5qZ6yEKGuXsJckdUD623dMC3/+bMFvON9HlJ7XFmU2H5AhuN4kIKoMC3hPtUpc
cb0MAlqny/F8KvxlbDyS+Y3FdCF2edtK2r3Ay0zUhX9HBB0SSOCMWUhNSFASyoo5
yEHdBF80qA/BfLkJzLvvw6n59OugKMDtt7VOtTxz+FcJUfOUCNR1rt7UxSd3EPI1
iUMkP5YYicxtKKLbg3z/1VbYwWk8IJsahlrpCRNsLoT0jKV1nua/KTsgLz9YJfpy
MjzyL9+3G3ewL0kn2ec0qfn9/dFF2NASvekzQX8h505xo8ZOUJom+pitshVkSAKt
vLHd1R7Kn+G8Mao96N0lBAR9dlwtY3C6XXIR37265NGo+SujYUTrHYaIFo6OUTOI
T8afp0x5jW/I8tvY34WkpjpbIG4xPr5LNtK+Kp1OSwG6sC3TO0k3j+MgHn4OIipz
bzI9yKI3+aenmeJK3HigGNg9Rw+82oovkF6eTelXGS1/VmuvcU1Qz8CeHpAOTOVH
WqdtCNya/LrCDPXEYu5h4ISlHxRRO5alGyUbL3hFh35Erd/ZDiKCG1+dWfxd2WPL
u3hD5+byrK3VFD5+mVW7vzFY8dYWsasJ2s4XgrmpICCZbVOWVRn0SBu+FATFOCfG
GgSMBmGn+jP4RBGd5bSuCCQgRbsZg5L7yPz+IIMk2bBHW31iw3pSowAb9/fnCG6K
JZI+S4lv7Ie3DGInqBVcp0FlPWhgWvvejU2+FFXzpO8THTBBegUKiEFCr0/h50FB
psakLt5rByx/r16JTJ1DhPoRLtA3ruglTMnsAcqd2AfFS0pF2YN8kGS09mzGbwmW
LHnzeVYh392b1RBSFBaQ1BYK/nibRKasQO5CpD+FcjDfAM9bViymX4ADPGKdO8EE
nvjYu66sKOqZ+KsNQud1qYaELiHv1LtNFyOknXfctR1vkypGjWJn28r/haaPI1Vz
pm6XWWuHz29j97EoDHVzXDITjA+hgUXRB3PkYHxkBN+JgSixuuSZI7gIHh61cU2C
NV6NvQ+marZDeRf/bDJAVrHdiJaep79ZkVhNuNHa9iz+tybTwJ9UHH2eODKwP+yl
r57m68Y3qOYsYqlXGaMZ1j+pM0D0+s0LlOH6QVsKU7vgS3sSRs1ufC6PjMjB5/v5
ICd5iH3H6/eXYlJgTlk1z+Q4eCV0C8qknUPnDNTTKlEgKJK0t++7+3zS0FVdqFAr
xO5uba97TZI6Wx2WE0Ted/yCm1XDtCfx0cIVM8pLqcfNUspROWum4hrvp0RF+4ul
nz4kIMvRqvojB7KtTBXjDFTBs/XdwPNBdYr+jBg3SeNGxFhVdcRItBIs6rgtPuZs
CtUJcOxlFiZFDbyf0Llbv0BNC2/dRIn3HHtTmg0EfD1W+G+4FDtbWW9Gmo1fKurw
dL4k4qJLgP6RMY6nAtpMsuOiYEyL98OEwH5IB5u3ODmV7yyF2KugROVhhMtq8TAD
bsLXKE1ByEtlc7z66VPDXU5gKXewCf05sEEFABXjVSEgvcTZxAKQj0HaPl0DUb5j
7LM/jzsPyxcl685Z2I8Wcfw55IirY3ev0p4r/WKyEiZ6rRtj3NN+bmqicZxE48jB
MZH2kz28QZkHxO+JVx98/O33DRTLyKnWWxhUBk3w6wH+amLKUm6R36VvE1TQijiw
wW4CmPFU+BpoZjmwhQKX7egzL1x4mYmQ7ujnnxwIBrgFGmWhrWhoDcoZdL1rNh5g
MIcMvOGzBM1X0i+ktm2Xmnb4st6rmItTXRpRsPsxR7zd4EInbGK+gGA0y3/dipnS
gw3VrD1I3w0gXR91Yb+ajo3lvIvxfVMF1VERshExsRUuUJ0KTVZONlDdqbZgHTKc
PtI5sjgKqFIU7bfDlnzYBPVzyGohS/7prydukHXOaz0qIOJ22yC9fEdnM9oemlt3
LZKGhqA3CqCHhRcLEW8jxHtLVHZxg3Bu+qC1G4WoHSNSas6irmcfZpEnW7i67q4G
Z6FhFFQv1HoBFUMchsJEHChaaKJfSmIDYuZUA1UU7gSTDvDiZ46EMwJs32ffZ8tY
WJAa5rhPpOW6+XSNParDyk+5YQhFlf2FHIrKHGpad68v42uSsHeW0/K+zakjShH0
KdlIkAZq868V06Ijmk6vceMUlSFpoQMS4C80QwY8ImFtpJ1D5Ar0fuIjZ9AqGrpD
xSI6tBJ9+Wd5Rx42u3cCre+6+YYPsXx7+RV6RVgwWjQcSW6jgZoCF8NYM+uXCrfr
WHZmxdrvuPMxEDF6pjiURVzuvhsdb+/eu/9SBc33WwTHdVYdwPV0F60+PDRrWMCX
WT1d1jsaBtz3TLaCMJyfuoMwkHMNxhJcTOirZ3UWTeb7j0+TIRsbRrd4DKEprFYy
xRlZqaFyFZOmaSUFLTmnzPdrW1WDTIQTaaNM5loCvtlKWJOXPEZ1KiO468UMv1wE
vPDsFd29P4CcWCBUapTc4xZ4fS1b3ruUsv1s4G4Au5vTP6slnpWWA36D6ePUd2GU
HqwjuG2Ma0WDMeeb9/zJk0Tm5QeQ0vZOJJKod39XlOuCV3zfimdcKOH50GfH6JYY
4/ZdZt/JmI9WsgD2jj6/IV/xwsqacXNYexNpNILlLeW8sRDDy0A2ZA7qpCS6A0c9
Xi8aP6hDw+puxmwYcOuqPCtQBrC/KIYrSsaoHUtzKY1H1pXMXvps7mpJneQ2BPr6
XXO+hImqhjBCjklBYBsDhYnmjsaz4E6THeI7z1ThJ00AFSmftXFVIxO0dS8MOENN
zNTSbm97eX0hnSDum9LcLj/kGHR0FefjYYBQ94TOwAkC1jjWiCbk5QQyJ07ptJp1
KcQWUqSR3/9odl4YbncNKP8cP+9hs/mKLmmR6RN6kkwPJx+uefPxtDiNykdkwWhG
bNk6O66qhDSDCbx91OZ6zKU/mYgEYfew5PnR7rVghDkxRgJdrUhFUV0aAN9ZKkqv
PHFce/ZrBO6jrh2EY7HVp7mK47+kveLqfx0f1ISGIHP/ARd9nmtfNTr+zcOTr+I+
/clFS/+O5SZnCPvmxJ7MiJnDYyStOSeRI+xhmtKvjryYNnRE3CTEDA/eK3v3p0YT
nIJr1cvCBj0fVLtTCPaMVrQrPTk+UvIBSgdYkykv5tT/lfYMDy2pXhAVckAtO6C+
xsiC3fkcrLnuUT2vGC9VQ1boMzbS3JQA5rf+66yffKc+fHeMLzbToR3Jk8LHWgSb
vMTAz5lpBe8sxO+5qY0UDW7TEpBmhtcpy6BoSXxmhac7epwFeM8nakusFKadl51z
kNoxxazjLr6ny9kUgk+eQcStpH2W15BhdOstNNuAwcc+trTCeyRKlnKyc3tn0olb
Nj61NDaEnCjyofEvA6Ry9AoV9XO6n74EkiAXBw+hrParDw3Csedl2QPFnnk/Wast
+Kt/nFchXgVN6se7Otuu/uXMR80LNl4HnGNNZyIJGgyhV2hWpIuENHQlv9he+Z4+
1/rUD7Dt3hY3tWLxDIUKH3OdV31/1rfplryeSfn+2C7g27yd+igDpemCLHf8+eNp
etZhyD069n41yUSjBhFPPxaNclyMGJI6CSrkYh9m8pUSEsRiv7IF29phBlZtG8/q
544DjB2QQAIMNKc5qBzsUWUVySjcTfKw+WMBXJwe2PlUBErLPjorrPEdksbwRFxG
37klYFTMVIHQvcYhjN/hTjJUHQunl4hvtZJC3ydslGQD2fEMNOb130VYr2jHHPTF
s5oFTT5pI7HXkujAkV8/9pvakADi5wGaU34QmOALfTOQXITiu852u0wHNQvrRpoQ
PjXpPFjMtomaRYUN1FHUuef1zj+eEfRDSH9rUGtKWH8eswHHDoBR25fwcd+/eoys
TMy07sKpULIQj4IQv6P1EFAjJGMVeyGBUVtvsb5V1hDzXZKwCoLhE5y2Q+H9NqeS
THPsGHpS1NYXcTFgEb32lvG3twF9yTla6j4NADrhdWJXKHBnt/OwcYj0hovBUfuz
EsgsIf1JXCg5gEudtSnRUR5f2rsTKfEKFRbti7BJSWhOMDIBOpZfJ7Se6RQJENl1
BEME0Sdu7aYJua4v0h2xPhX+ZzOKA9H+Npy0TOy/aLkrn5271FO+vOjvERhFQgFl
FwcbV3M96z46p84eupTsT//8Ww7BcgyO0zeqwnEQgbQFg6oH7z/0mDyTdP8i9Z41
hWgwPG1e7Bh+1il3HmJL5SzHnJ5/B8Ip5vnUPLGsalPryN/KUdn773IoqVDZmfL6
LXh5cRQJxSVszL6Ijj9ny1F1d6RICg255JsuVFLLz7SnUfwUzA+IogA2vUHjc3f5
MVfSH985by0ocMDUe0C/xIZW3NT+y8SV0hcxFZI3TzbpMGmk/fVil64odVoEdJfP
N4p7VJF04OlcsVwyVXu2T3hnSbbafNggNOWbFn0ON/Sq1LFlLVl4oSg1UO371ddo
D7fl/k3kDHsRp3WMQBGJqi4CeR9MVMm2ufgpGDGFrMYQOmzm7KWN9NGu/vqfTZgl
FkdOLtdku8jU1LZ9//1Uruy/qASIZfjxEeGpvHGb2ZVZwZH5eyWC7/eVwj5N7gzh
VdyLtVKAeXeMTs10uVe3nt0PhB7AEBqysgvDY7n3V7qt00EoO7vrEKF4EhDusdG0
y5PdYkY3C/i+i0TdURbvFp3OSLQpdD5VrRtdtyD3GnXligCc4P8MWixt9GyOJ4Rw
Ci1HwMO5mBQev+K0+21GoRowcHeVkOMWrT9cQ8jkpBzpmekjv1yJNsrpTKq52qfa
1Ot0hdkUGOOqUWT5PXFCRrq91bDBaPzpp0J+JljSllJFsOaa4eLrLmy9zoWUAsMO
0X+B2VN/MCltig+NHr4JZTEub0YxpzInVZ7ctfNDPnUNWShUY9eOBJfxAprNaMSj
JybyVlSrQiD+aMpDr/9OpeWDOZMWcG9TuYW1+xIkmN1HL0iJwriXNEqFZwoApTSO
uX/8Pv6E5DHAobwNy8V6KsyC5GCtMxBehdO7En/rKeiyUlLB+0fKE8VKpVmmKrJL
VIN8rsipqA43+KOKHIbiVNqkUTTklRBRlqxYgQ1W0K/YAQAprWyMvJ3qCwTuhCUJ
VWbq/yF9IADRrVyCe8GRQaclFU4IT9afSagWRY9VymvkRdhcy54esgDJ5pSTSig2
O2NYWPMzUreDpU54UrY4KQgEUtnhYTAUOX0kX5bNnvSrgLObkd5oCMs6DeM2//rt
WpqVjs5u/SV9Iybfc+3mOL5P0zoIq35DHKBsrj61F/htCXBewVinRKjfhjl7MLKI
9/Tk1otjgda8/ekqNzpdqqlFBI6F7rJHHUMVG0zaP9FOKIsOLR14fym0gAFb/oKs
ujA5dF6LvCM9TcmL0gCWxo8wlEGujT1vc1F3orhyu7RnjZHI5xYt+W1w8pLKSiFc
PIHRIM3HoxUc8uH6fYCVSkz14cbY1rauFACr+pcw8ZO6rf2QlHhEy+ChTSmFsHQI
VI3vaq/BDZAeT4EKxoozQIJgfN/VNDmkc0UZEj5aCsz9v5UT7AR6sKrStZxseLbq
gBKx8Qku5IGvEe5D5//vPjbWtSxDdlvHCECGf6b2bI1Sm8AyjYeKRr8PcNj1AADC
2K52RM9wFikg64YKp2y0FXscmCp7HnFEXpZ5ygvjl0jFe70z/7KQviUm/pweE623
kOf61ugkg2CzMMGUPyQTJqrKAkDx3fAsks81SLNCXD6pTc4o68V7ru/XMxUZYJg5
cJUUtgfCa+E/d+Ud+/aaaxmxDJhexbYOeZVu7OBF3PASUffhHZyQwm0qXPg1FlAp
L7QGSct2yE0uDD0ov3OorElCZm96cFd1G2hR1XT+D4KBW80GG5cHzjjjxVABjp1l
oNtANOKDnfe1RP9uqGgMyPpkxm6jn+fqCl4FelNZ3bkvi06D7cj+2ocn7NZnzs5u
1uhX2qC+Xrwt9bWZGuTQhCpxNVNQ2jjHBh5c/WpEWBEn9hvx3JF1R2TeKQz0AZVi
eDrHbgbV08BqQtq33Z10H4qowAh7DDWfeKc2LzEapMzMwLPS3eoXCmf/+VoEwrHs
qfr5L7ofJOu3gNKgVXJ2PUajTPErnDR6DW8GjiNvc2gVrF5E3oJOreiPx8vzK3wu
RH9yik87fZK+Krj0VRnvDSeqmJBLmFxUnaDxr0NVB3b7Id13HaMDcb+6fftyeYV2
loOWh/g6//iMFkaWO9xkCN/BFjPAFv77iVKQ35xNwdJ2Vq2SLmlnUCbsQ3LLPdSN
IWOD9MaXxKOGv9oYKrMGTyUgLp2WVFkcTf3cmphbvqjkZj6q3JB4dtNSvOoZN6ZW
l3RxOVpdDh0TyhrkdBR6Z4mQjQmCx3hyRGldqnADeiMvp1O8UdGnwTOkaA8e3DaK
KwKjM9zPBJq74zGwc+ohNz8AO/34JlYPhNiV1CCNMOknrkG80epHU30QF46ajmkn
FyorLnvQSNKxUPRRvDWeuNSHrAuwC/IW6AYzAMLB1n2uOotNN2BHj6/47RSKuWhy
SI4sbU+V8aFcuZ8Axw5YrlikncQlApv58+FGQfz9xXK9PcCFNRvk92KUeYFNOHXI
dggA8hf6RYHdtpxMqVU68mSanljQ0mQjLl6chAE/IKMb8S1f3aY91s+Dckl1Prtp
NJf/EYRTdOS5ovP9JF0TG9OvH8Ctx5a/FJo76svZJZS97yvuw+82Cx1XMNoYNJOF
VP5KY/UC+iY1ZxW2bbHquvHmqaekwG5e/X3ao2xCUYvkjv6GFT/+WN3WeF2kfvkc
iW7ERXZsLMix2TN4YXg3SQl0z6qv98gxTmUNcZuEXPfUnROaN3IFq8i3afmm9xGO
LJuhdEKUpK+C7h5g8JYM/u1ger0q9lkwS3cHa1O1+H0OMi9rl6z5/uf91duztP2v
D/nBurcPzibLYzioaH6YhNhHpd2eTzrPI4wWZxz730NB+9Ozbs4ZaIdbEuMWaNVl
gOPmNqxjvGqxUPOlVh0F/fW8T3/SDmkgBU/sEmvMf47FzHFfl93dsTG7FtxbhIDm
I+oVCCwtdomF/kF7ZiBC9Rlo3hMEm3dFEr4eiBZH5J2kNY6B7glYpn5H1Tpv5BCA
a5wBc8U+y7cMukRNRGpkbM95VMKmsu6P/6+wpNMaBSWdbbmFjvDHfdtzD46gKGZh
wLVFUNXIh7zeW5EZqaTd6h9BCv1iffSkzpG0cbO4lLRP76rTD+UNlb9uo0Zrhf4Q
X7dFqtkKSX3r1ZpuB3Y0F/qSDD1179+PrF56uH6O6iASlagAcA5Jgbe0SHV3i6oR
wDqin7rEHLt2MlvUl4leUIBe9Zd9NlkDytmbOL+DyZtD4N4G+FMXXHOvVP86aZVw
6sWtA8pWjhkkTFT8TGiJRsx1jF1qe4yfUxO86lDYg6sAwyFAbL7lT6b1dYrySAbR
od1zarOOiV8Fe2DfO0SuWFw3wxlnZZLiKuimGlJpgWi7CYfD/xSLIpts8FhgDuet
j6T1Bwh0lXSAt140nhfxsP+Q6busZ7K2aycQAWtoGPxfdJf6je0rJxCY2rDTTbY9
IrYxUcmtikLErh9UVJCRyBVf/Z3UIvx+2syOECv2PS5vxho1B2ljHrb0WqPxNmQJ
7L0Wtctu/qTFeIaRbxQ1luglo98IjmwIhAIRgFKhdEesbfV0HOgwXPO2LohCo6Rh
9BoNGBh8znnD32FV85SY9Hc4kIgTpmFJQO9xvnNkQ+E5Xv6iRr+N+1tnsiicNVet
w54P8KBHN7t5RfJ0gxZZ2S72d+zipKi4lUNusnCIu7u605zErQzET9XJ6KK0InMN
iWHFf5yPVIfBTsyD8GnbD2Rj593VuPfu7vX+MSh0NIEH0AIzqV97c+kwuluSZb3z
1yc/6uD+ygGtG2xG+h3SXpNC/D87kc3et/1d5bgVObsU5GwOHxEBfhRNrVFSjJgX
egiqCVh1h9D+UIM+4jlciQQi4jjZpgiMaSLA98sWhNy+WdRhwpaz7Cm3UThZm4U4
HR5jtHLm8ioVh4Wl1kq253WsoVAyfNCCDIzqbNjBWK8fpLzS7dOfwcLkXwaiM9NI
LehGh8+UvmaFmifr89pb9oZldOAnXRJyycyGyq65gxUsek6/tKdAb5vi7NG34NzL
nUE9axh84KF7zuGwc5n67HZg7j+sj+ef0a/GNxSLlvUear8X1ldTJKbqu/xTDbaM
nYUe01IYCRtPk4Dm6e5Na1yhyT4zByC2DbuvD20BpvDdIMHE8V7u3tZi7z0rHYxC
pPKbAA09PhhshAxstIKstmsom0jmk5ukjhoJnIqPL1BhzqzTniJMqLLylm/FGKDY
kMmjqSNS2Mum3eDB/eCN42Ay9MI77stQbO5B+1ohKtXz2czWmW2MUN+oE9YwBbOS
/XBWLUcRoNXjGk8sE+SrTyk1ZOiyIcokvGtwl8pTtTdWvFTNpZpGINBSqYtybWQU
BBdn3+YDRLF7lkwpO4/52fnMkC3SwhZzcOYib6t9THSKDgH4rZFIrKoCLtZDB0U+
AfTk+4lPjzLSEr621j6fGlDKu8c/zNyMsW0BE0gh1LsryUL8Z3gn8p0UUSPB1PwP
tvZFzMg++0Bt1nZ90mxw2lmhP6PVrw71/Jl0S9ZxpzWrnbVVzgMytQjpKEKJ/eCq
heCKI4oLPe89nmdOa/9aLUmPgIb7tVN2eW6rNwHoYpYLozkVihkx/RjYwRnTlK9V
+osDP+zpSYxfWxCbNJpyUaQaheYlqoMOnuRhR6woOP/dRsQjkD//wbuVg5/zEh5Z
C1SAwdIHtSm7tuirNjnYs9NlENt02VM10/d1EyNApmZltiJkW3vRY7X2WjrwMaum
5cxZ9mHSiI3cTYUCMj8KX+3vne+Sxdo3W4GK3LMOnk8KoRPrll/LdYvedcs/HIp+
VGNzk4wiQJMt+L15fcDq2q7zksLUZLzNnZnDvjUHq0hiBzQ1XHJeWV0vP/6uUXdi
yv4ps4irWR13YVNT67IdIftxr/ec0leg1mTZezKcOCOnW1Yj/Dbmj78S4IafWk2n
z+WgUjLVO1VfhMhWVnKo3oC0n6HWxuN0qjVMsObRaqZbxfs6f/lcTZw4KUZXI7wV
quOA0Yc3iXLD3QqY6DQ9uMQc/WS7VNaB0nlaHUJMVRKEAPidDqVefCpqxY/In/Lb
VtPWu1EFTyeLvcRfwCOEMCI92R/cunJ1Tg8vF8faPTnU2pLdrmQhjcieM4J6O+MH
POlVesjI0fdvWPG6dWQukuLPyIHkKjhhhhcQf712VXrEgR4rV3QsQtWDi8m6O2i9
pfP0YMcHZWN7+cmgq/FIulKPAw1Q9LN8UHJf9z6L+edRG4d2Ayn/nD8U76cLPyjI
uLoj8jzJMBrXKTGj3SNnH+Wk4+OYzJhfRH0KoUhXuSda3J6WdPqmiNHUGc7g3Luw
UXmmxR3GAWogQWdKDSGWMSREa4HuguWLwfAKRKzMZE+1GVkRSYd9Lu2n/JUcOIbv
g/BsCqtihjZlfNPu7g22J25Cwh5IU+TnENiHadJO9sLZtMSsAJbFa85JWZXZwfuR
coOsQHAPy9EWTonHQotrRMYOLKFYUQvEfOnX/M/+HIo6iUHvWxtaQQGMBkPXaoMK
TmVU/q9EgbiR0OoE/YS11y7OHwsLN7+z9Flws0LUWWmNVrlXMpixLmCgD4qp+DJc
oZvnRJIjioAIkmXLeFCAOUQZqvs9LDbxPqLld6wZNBgYUG704iUxRWPiI/m3YAAg
dCZoiPJxYNk4hzi2tNFOoOh29P+Vd9MrUL9L2+HTi/lQgys3/AUuERxIR5vBsypW
gEoqd0uP83mmG3pwo7ttmFgAu15AnruH5UnKuJO8vXLCTrZugig7My1nLVc+MXem
021vOfsHT8Z4bgOhBHJDWtBqXFPpviHaF9pmZ47CKihbfx5MoBQTq+twXmu5ARNV
F9kWUf9Afkv7GFNsygN0WLnIW+4ugzFV9Uu53Y5KquVmCATtsBhIBfystn/eV0vI
01XOSDuxsVH268s0gNftrVlA02Z4hJfoYn4v+fSii9K13zngC9ZfSjq6A92kKfnX
0nlPXR5WCF8PHlCJ3jkgZRPLvgMTbcmCXb6cTm4LIdtZnMe9PirVsRZh0eynh1rY
ViTt0P/UbzZxhlru2y1Jr031aewqA2YqQChG6zDUI0bl1FWG2kigc2kinKrjt3Im
eB7U2XUG9fdgAjJ7zkWwnMp2bBa8sFGvUAQeJLXLpTr/NBZyPegFT5mz7leQ3vi7
dBToQL45KdtQYaSr8oJJVts0kbpj7bQ/SrgVks0Vrde6fvVWhGXWMHNI9m4JOBmj
gdWJI4SMWsrw/M+pTujpqZcMoPUzzN41JStbLgpEObswCK5F4g2xRkhv9YRiwTgc
aigIYSgstZNa66hbFX/NxHI9kGWvgQOhU0Lq1FZeZWRJDddTXzWiQ+M/mjeU/zDc
3ZEUjK+tbSZ5Ib95ReEXco7B0GmGwEudFMhKXi7huo/yb9T9hXihHEaNLLazZu8M
grMGN9Y7hr9I+KfA0Y96xtvlOwKbq+8lwLqUrUcrYFHmdqNnnq68WWO1T/uo4P2r
dOxU/TchKJlw8X+Xxnflm1wXvvTtsu9U1gJHUHm3jxoHMZQDc5TPp42JTPyIr7Qa
26WdbJfdYL/I6YQnwQxlo/V4f5WFpkNefxYKqzJe2+d/MuMzBEtbplcd7dxSh6K5
cru2YyGpIjaoNgarHIQByQ5xJZFiplU8IfzId9pAJw2T+lCvKeY/rBAfOXdo2SRn
jbyKSHgaUwAg9LpsP5gJY7gHQTfGvfogEgYN9uGmnCzTNeXAyW42bBRkJFEfhf0b
+DPuownetVhfuZ0FOX4/SPrmVF/6zyjUhkAcMFvPvYUWfWvJn2uosO7xKK+DlUpr
mLVoeMqQ1nVyP/1IN35pBqmaNpXg2XSxpBJasIKil8ZhMRW407dU60SL9eEx1m+B
PW8hUMimGvWg1GplTs4BjOIJXj4TMol8nT42jxfU9UPe9NBlQk8//jMc83uaGM8o
eRxK2vjPwJDoQW1La/G/wh20RYxTsfASAWXVqJSs+sB791TBq4H998P2fr9OKyjo
mcxwt9B59uGmYwiUpnG3ybNlVxxrDfEznJExLxdPr428QoV1uCABTDd2FulegC46
aaFNWpWC1u0D99xFKOsQF9sXAom7+36yXVIWz3m49iCUv62J83Km8XV8A2YLQfBb
f1rn6rfP+GO/U8/LpN2mgitnBrvj1sJbCWantXPWJkrgtFJzld01AvFbyfSEZU2Z
gdO6gDWud/JeRIAs9icJ35qcGUtSTtk02CukmbQG5FV81eo9chZbePPaZpVTIOyB
vymHT3t0bNauL2+eDItDK6Q9dGEqlz4QkdUKPHlCZ+ha4epsz0gg7rfEgKwYC46p
6RfQ8OpIzkrvpfOYIpGXywVPqABjJSt41LRjBMDG3E7lFuI6X9SjwVGFe5veJma/
2u51O/9oMVAzFedpIciCWVvQjFxRYRS/w3IQLwkyGVjGSNXVE+bB1H3QjSoho1pe
CJ8U/YGWTQKXfmg9M3SzGtcFXFC+UHq/51jW7BFAR7mZ0LRh9ToprRaQBgTBRg7j
/WNWdKW5zp8gX1rYpeOGRfadSXAcen48F9FpJDLgrNHTF1DpSL3SBHXUxanE0rkx
Pcd6XwDb7SCajlkMQIvou1pYOVBJrBK1UqPg3sw2JPUeZD0ZJXNzZxFZC5XJBbi6
DNzNe127mxIiuTu+GGuS4kAotfSTfP9U8EZjzq3qjJVCETwXziOO5DKGRwkPNweJ
q9fW2H+nNovpWTCwQVU1LwISm+PYiopjLltg0Ut4QhdUABGU0rayWFshV2yF3tyF
aX0aIuGfxTcYnqv3QK6tt3Tb9QJEcgbbPUsWwjrx4Nzc5gZtB+ELsuw1DCq1ja2G
zxFjq+kig02Ls8wDR3eu+awht7GfU0pdhqUl1n28KqkQHdYuChilRYIonvJnO1lh
t7vI6CnbCBB+6BJO4ocBQChX+ocOasJMCNaB3ZuPyD/4aM0+BzfuZokF1mr5waAo
F5NtUfyJwkyV3y182ZNJPrl5Ua2MU18u/rmUegPxIPaVASInG6wG3ruKEV5Fwj+c
JGZwtkVHT3+L4kYBOudMkm7Oy2x9Do3ruHpotUwPqAjWUFFSjpXkhNVM5TPYtsVN
qKpQZrcr7CjJ7lrrrddGfhrjCs4QqZGMcwHbqH8/jGP5twZ/aeIihLbwUsj5fvgq
DB3JqIuBpIWSh775orfHxMtaKYfvbjti/ibgSbUqirBiDpwwHTfBLAY+Guqwvfak
ZWVX2/m4UiooEaSPtcMFa/rOxvJfnX+3EztmBApS0oib0fW1nkR3vCnj5xEJp/w5
uMXNCWJ9XoEZVMbVIh4d2ZwjQpmHaENH1HznQK81bCSCqK6yRXyyU432HQuTTAO4
t8Cgu/4KFmdGLr275dg4QWQ/eOcJA/qTAteeYRxUAii9bELzomeSvJ5jwMXhRPGV
19kAEj3JQ6ikMulaObQ8sFMMqt0y8+CILn0BEu94aYVEL7DgmkVRs7E0s8DnbSDc
bzCuEYs6uyAWOzu0yz+OeIhlqVSDAoLb+sVEfRqzr7zRM/ipD67Hiy1HHV1Hzqav
L5aqzFLGnFj4jNxfAOHoEjOWg6YmwvYOpLVWWTgXI0F+y4+aug2jRoJrVuhEIMif
Tz+XQSouWL5tN5hk4/85ZU5f/l4n594G/83RGXUgbvB0KcSQS3N30UAsHK9Lbq+u
LJC0XyFLyP9Vt7WCQqpSNX15vy5ucGVyFI3yAI07Sk+kbSxbp1tI3JYXWLMha8eu
h5pdRg99dkiOAcy1iEKD/dJ/qmkwPR7d3CXWDr9yPWnM0DLkaAw/T/qVKUnaodBs
4Kj7wz3m6YEyvtyU/b8N3Ra/YlQjapm8buZZ4XNp+sp4Tr9/GlTyXTf9qhbJ0K06
+vBV1hRS5SRS20tUAPzEQH1JSC6rCq1U4qVRXsq6i9tC9aDcUJoXeMb9fTioNxUv
4I+xQmsQe5v5X/+E6a0cJVG6CX1tmrw3dZ4PrPy7rgK6AyznNcwupocpsUouVrEt
3qoLQoiIPQUQzcqFOR6TJikpua3e/HmtuUO40o9zdSFtyT7oHs731OATEs+AxiIF
xmpiHozr+i25k7IAAqsTaUTdtPfbWfTkZcKjUk+sStcjpgQO3KkcOAh7BOIpkL7L
1803sTNituxTrBpT2P0M6un2cD7/hOYRrD+YVQYr3TI5lrzNsa/vu5d3xoOdeEw/
O3CFL9/Db71tPkfs6Q3LlHzzsEOcCBZexes/v12bbRJNeOfYBitea1SmGoieDR8d
0zI/gad/tOFSW949k4XVPJQkzE1rYNPY2QVbg1w2+G7DSqx2hFyDLBvkIt58WfRV
IfRXoK0/rmGqakEgn86rOvyQRLiPjYfrhvWQma1/d/vjJHH9t06gK7YUjeOvYyCr
39az89kKQ9OFtmpShKg3SlI1HGCplLQ1Kjmn3xPbXdr3gQ7IzBAAXF8F9HD41/5G
jWz1hCvKo7tfgwGY1AqNcU1MTRl2MnyM/uB02vBquQjKecytNIr63yUd1kjOLtr2
+gEzsfpEGX+SSfPWwLb+Uwr+df5egWwqFrPkZ0ObxE5cbwdVq+cQBcZN/riEKKzY
ri7loDFGO+U74L1WMXxpknSbq+LJoioWV/RzRKnu6xFburFuuor/bDkvcpZ6cqj8
rWC8Uy+emMNeYCxJEoTsOfkwICEJzlqOoLFqBW8DiaYqjwWprl+faqrOqFA1/o77
zmvEvAtXq9cIJeGimbETmqb7Ql1MwxoBpNQ0Xg0m8lZj3piEtnJZ/WCikISUrM/3
7oquKUT5ULxFBMJ/QWAwuzi84F27Gh9tx/MDSQQQp4weplvINrVaeCh6Izy3GVpr
91d07b/7o6I9/cRTotSZHsdLocZnKh64m9oo1WMJbiv1xX3GRubDZSU+rqARsKZT
U6gStm7YQYA00/EjiWM6iZxdUdH9LmM+bIU/57rSd0uvJaz309uu/3A4Lr2a+1x4
aMAeZrIoWPItfRRVXJFz2zg9cesCwChO7QowWO4TN+K7JUe3fgq4jhKBePN28FOV
+2CgC2vj1HXnUn1S3fNQFmnyNYXgN1jKxc67DSrgh/apw2w6E3U/FxPQYHhgP9tc
EQqCY96zU1wGllE/NsIj6Hc7N3djJ59x3Vt/YEzFc36T4IjBICC0aDde+Qpea/3K
traiE9Vzvg/iSXH1pSlvhPs6Ku+juhNzyhgyzBTORa8CUYUORqDSgGw1d3Lh+kVG
yWANj4O84v0jviaeZftEWnHupRMecyBnIccBCNey5pdiJcno/bvTQE1WIJRjtxat
QyVsDm+0ixyLDpO/KRTO7+L8H0dHL/FaCs3dWV3CP6bQUUfplt1yp8EM8Ud62KLr
yErkx5J3Mv9xXB8pTA4BD34rulCtjjwKLPgqEQM7P46hkvjOwtrE0mmzDzEEDZyP
TYhpfEDmCEOfKLwoDePRFYA/sOFZZncdN44G2a1SpnbJ5P5o9EQIC096mt7xBxh9
x+a3cuPLuVMzwjkK4ZN2p0fauksmFwHTEfhcfqK9hqh1RrwcKz2BY5ycAmQDJASv
m9PR7QqsFbHxPvkdmO5s1smd1Wp86rjfR1i8R7g/IJrEAAiFI5iTXhhTXgYpJE0r
M7jqwUSKAVG3CUpZJFQ3bsfZdoGwqDT9JZKgUauunDLgqaiy6CHSG8zZbGyxsnqd
ScrSUd6Uhvj692Osrl7V5JPHq7kF2TNtH04fnCrOwFgMadtcw0Mp3IcY7RYyFkUA
rNSpYa7eAxCKE7N+tU3ZbdJOhjg9dF3+DOg6CKDE8zsDUankcfzXU0I3xEyYPIPg
1pU9GaetXX0/8zFhZ85qNfZSj7kTENzy5nRPfYlhjnsMbJtL9AHH5B6zWi55BRIX
Ei/qrbjNprVlf6zkemZrN+1j2g8I+8zrg2byBbGKJAf9kDABY3j1OzP3CobvyjN9
SmPmx64GZrncTeY+b2fMJdknT2KPuBEJxIMBm4VC/4bPC8MYVJEIjq/inVEG+f+9
lxshpH2ebXqQGeA8JBAHPobsgquTFI7V+3swlNUT32sl+4Far8I5Yv/pg0JQECd4
J7x5L0PpRTCPs5PuD+sMZ/xJsX2LI/YCs7TY78o9C4TQq0PGznxUQXnrh3QOWVBE
I9R4yVaiYvLfJc32eio9riyFYO/3O6l6bX5UxBwn4K4DrXOIEn2DfnjdiGePVZM9
x6ojc89++56IKPjq9LJiE1OnZGtYWpb7PoRi+XFrKAPyY1kAQaw5gGGOYhusARFl
dCHSMkQ7N6gd7BeHhEH6te+z+w6QlIwbgBQSpLbfJQa62NPegg5EXyZk5kBgEq3K
qcAUkYfop5sUthvSrTpUlYGXzhBK6kNuMG6VHwuwge2Db8RmLrsKpDvE3XhndAPE
c9LT3mCAWwgVVFVwe7bPov4UTxQWxCaJvaaaJuk3JqIWRVWwODjsdhs2Yv5+kTgV
NCdNHQMlinL/+5PuMiCSxfgQ7CjJ8wHtGCGoSBqgFOkP1AGHTp3/jGtQ9Fzc/LWJ
KtpfhKPAXKSyoEcYkDQpuUcmpkYl/d9VtQk0yJS+Jj3mUE0116kvHulbXWhY08uK
i0qbJ4fuqm2oWDx04faX2/NvVe12kq+cO5xsTG0xhhBXdyBoPM7e/WhkoEx5oQZM
c+fIjbDSnsTQ2PjIwurzsNygmiOx34rUKLsO/GT6NUlW4qBv7wF5Cx3jxsTVSyi6
0jULyXPST+MOSRZB0T/OO9OlcSrdQTwYR9tzTjBiXMEEpLLiNNqnExQ0Fxf2IswL
bT2vaZeOsDgnwXunNSqdSqrM7cZsiGM+1ty0SJBnV+CA8AOODHAHDCtkymh1DWqy
tlOefQIPV3gVoNLUC1xOmLsALANIQBC+apQVeMHVkeYV2ozdjffobhXEAGgbuiB6
eM1yQesmncLSZA1axNw1+8NxrZYmGJd9kj5R0dTzO2u/j8DxmGxNnGJLFAgkw4d0
0pXAhTw7Ay+fA6mNWMm0pwjHwruT5ULZ1qXhZkrIfBBVvW4x0RCpuJXDE5ZlA8hy
OSg2dO5JaHaLn+9hWhcTzzhiJMrK6/eEqXdhnKITPBjad4Ix4r1HAqK1279mr0/Z
h4ALVCrO/SCnh01Cf1J1f1lfEPGnZMhGAbt07z+81//TlfhiLDtOhUY1Sy+CjMDC
zi9YPQ6ddF497twe9NzLYZbgmw4/WEpu2tJtu/BDkEe40fJRJGEp5kOid3BOue2Z
SfCQhh7D0oHFZ7kEzqpVAMJ1EDobwDrLFSA3ibnYM7KvVYuldFh4nwQV5nSN1H0H
saBEr4TN299rL9m4eiBbLptDfRepyt7Ep5hjLmy7YqjQBXeGC6BMeQTIeIEyfo7y
abZCjm01MoM3OBYp7N5L2xIM3nELDyte/BLqX+kZIJ0ihiKsX6pbBEMoHzoVd+LY
0G7/r+H512tPhdHTlJFqMJ3bSaET12WgozGw7tzjojiWvogarn/unhFGdM2wW5e2
3K/srdsWxv6IxYjcrLzqMnkFLSrReuo/bBm7l0GJ5+HaVdeai+p9OQnW1IO+kVrH
LR8frlwlg3xz/fw7KMiO5WUSFe4/f9DxmFBXH/1LG17F9l3NgzDVeKg0N9RQzvYR
LPnMF+fuUQzz45flbN+sy2t+PbNYuJbMPl0UYAle9e8xZ/+hG+auigN5RwcrnLdx
JkaBY6MGOorN8XL/8H1Oi1xm99fZCWf219QcqYdnVGM9x6CON4NEuo81H9M6um00
Hqd4l+hzOci8YYO09ftEnldCdbn9qAyTJqUYnPXFSEEo/Xl6IMRPvNgVNX6qvN7A
A3ukSFdCLo5mw0BMRppM+q8xLwGr1QmU99THbxhFhi+ETm618IB9faLZdebgSbnY
0RolOoIQJvHBpehRq+U/DDS9APxOHSRLrjDwewQz5StgP+pgE212VpjN2k5XIEzq
DwrZWFi+bNMr6Xo5V23iHUDhKIuvFvhdtVfTF46nvZ6HpVL4VSPjfKcppHqXBRKU
UUy39VaorXsLd/wMd28mZe/1LfrqEJBRZcvUSbG0J8fI8RLtEMaRfAX0kke3xxbF
BW0cpS5eNihl7rsimkWpCOkkF+mO733vV5mttTPFVv9aQJoBA3CpSXM4YM/JkpRk
6v9q7YjmWt7b8Sl2B5fO9xeTFSOpoLZV+QolLp57cKkutdfqvRUOo8rMyrJZsJ7Q
Haoojdz7tBOQp0z3hZ39Rn9Qb0jywERhholhGsYB+hspUKtNEfGYXMlqbo9GoxPr
AJrDdORsXNkGYUtzRpXGw+IxV0cYJnAYq3M/a4+Fw2Z7ghZ05Q5gmGCU7Eu7DUMx
GwE6sO3UIQcEtx2W7Pr2bR+biCf3s2VCA6PeYj7qB+6OBrxUWnc6xRD5MgBSWomU
5giKYBqsLQNlcqiu3xMyzpD9r+Na7I4HUHuXF/Kjqs1KvuERTSIrYPbLMzpv9Z88
46wJX62kucgrtrkHpPafrWmFzdAbFPGreWurhFADBjaKwZXSRtDMeiCjuKt777B+
4CXW0xFIbXRcd/peRbuQ/33w7d89qiSFktMR2MLW8B44w3v5Gx5dz8gywWqRyK24
fN4ojJnK8NhG3fOr6Zn0y5dGjjQAronod8JDuDieC94Xy4KZzYGSbXX4FAiwiNIH
TMtR6IoiqOFGEmFaKpbOghq3AGCCpvQOXqEE+cpqp+0Z76zLtDvihA3dObAVVwXg
VD/93dhCy3HCX0rLB95hNgv2FYWPBk8TQOqGf2auAGdcGd7lNMwgoQoQcFRYNX3+
cOdHUIFeDUDBcbK3Ft1I0Fv8t3DQcF0ZHREfSn+K40T8JwvgttkUt2ZqvtlPmI0x
uaO4s6fJwFtoEOw8ysuX6GFsTmkKartWQK4ocAIyzOIcL/IWhYLqf7pLs61BgY0A
aEwfF0kwOkFkfPXYkLAPEHy6lhm0gYgoJ+x5r68/lsrFdkV6asuW798424UFBG/O
ifbUNWdHxzq86wG5u46P2cM4fClfA3ZF25QnZQqNhHm7vRUeWIe8rRtJEnvjqkf5
arqRAJjXuwEK/fAUXhx4qqDEplwFH/z7KDmpaoLsqzPKlBuvTqxUeOuWzPPGWWk0
tTsV/IAwR9IMKntt6tg67/j+/PlRJQs16BUE2C6chPXZRVpEeWJ3UwV0ImkuNW7N
PEJPCzlj7A3AWRqewVBQ86AUg0bp6fhNUuZKf1YSd4dcqR6UWdn4fNe+o2jPhvZR
ixV8y/3rEmFVm67dB7P4V7ZHCvfQF8inogVGp3w7dbvEsrj5Z4O72dERWChleiAV
obSFduyEt8iX14lHajqgtK1BijVPzd9UHnG/y1ET68sxheXj4oFN3jg0jlyK/VsZ
egYWyaoeSxndZ0JMDZB5/bI7ztfPNgJez6+Uix6YCk9xEug9d/WmbYVAwK+nF5TH
Uinnu2XNiffCafnTz9XkBrkvW+m/YvyTAEXQYb+4v0aCEZaayZ6w0f1d087LIcWy
Oi4OUpUbYvYlVKZ+Y0rq3DYPw0LSTq+rQexDKzvklOveldufGs1TBfIFrn8EMYJE
QGboVNVHXfrf+j6rrH8G1G3wFaZcV5JOi1sOEC005bz7VPxDFWKcdZr5UKin4JGL
hrjAmuUM2ijElb2q+25lhVZMCPeHp5DGMKXXR5HEYU1gnwp143WmKEeCGH3ObkA/
ZQ0Ub4gvdid16GBXlJjcI2xkPbKo84RCaXqcGmeDJgUvI1SMBqiqNP4DxCGSzf6u
x/nYTzWZmgiZsdR+2BYKHMnRqeFKPG5HukbxdABNywTwJdUlEfadc+u8zOTeyPHP
f5i1a80S+9JjJhcIcIlzsGOsQk404706cOmI7Iq31a7DmPGmEEuH+YFNKS1KWkau
N57WHja/SmbldIaTJKsJ30PASw4UhuHsK7OXseN4FnL+ZQ64vNgsl0rAfLDBaaHD
z4M3x+XyGYYyMBmi75YlMm5/XMX6Ta7pZ269oTcO0dQQoj95gyXdTHhvpZuhi32b
rSjbMB5WMyujxoZ6EkS3IHxOWWChtKfW4w5d2LezLtvyovBVtplrxXvrSfTAPAM2
BE2bNjQItHj7L4CTScma1HI+NJf3Ufpp2gbjDY9ECZ7DNZVvu8KJhhzkPG8wWm9b
JZNfv+Y+jhy3R6OvNIPbV3CyJZJyLZGGaOw/0DErEfiYE16jCgZLAHSVyRG+9BsA
axVCtKSNo5zmv39bXr/JyVNMjRS5p36L9cLYqdCBMeoPwWat/N9Q6AqGYTuw/H+c
UjAQ50qacRceAkAcow0q2KvGI7vF02iK1/p0PcwQaveIzfPf6oSd21IYOS4OiXJ/
zMVpni9QbyZbMidUwcHQp5A2JDD6F5odguR2y6BsU+LEvpgLwZj6RTFZB55g2zcp
q2tMAY0vr3ygwyucSELTNIqeROck8lsrXfM1U0GWRVU3Ry3lRKvjmKmZXuJ1CPPr
NltMFkeq+bDZim3DFI2LN06ODqXx5uOb2WDwJSU7Lq6Be4Hij8AdzP5aF+AXpH+j
QZSg9PXo6uZW4HK11OqQLEHgNWbujzfbXWTFFSqaUuHPa0t3Ad0WeZYiNNH0yRKt
QtHSzRawpRMmpWErtEtNwHX3AX7XCGloGkXPs3menXfmvWZG9ku2wVUX9EB0JYwD
YbOvbUc4x4IHPw++rm3+Eef5wE7p8KM53+Pmbwml4f48OEySO/7O3rFx2H/ahpAd
0abWHdtj9gD2eWnwIUXqAnGiJSc2oOrU5FUj8xmmh6sfNSbRR79MdrEtfxnikxuH
QeFTbmClL8Su5qDoPfLxeUq9KC6WaoAKiiGWPWG9/IuzEsrtlOP2R2OGrC9ZgeFC
lunPoFMWtces3d3y3unJfUeazLltjoZb07h6LoUbGzxQNgfJx8LqWZkKNJzp/m7S
ee7WAFnFWPEP4bG2EXT4uPFj0pT/1mMYP4aHbl5pBUP/3g4w2G7nnQJMr6qYY683
sS62//yr+MVTnRWRbMT1UDcujvTTc1DFzTrWJJDr+0Pc5lwPMEUHxnVCdj56ULFd
wImMaevWgn/wq/qTPZz+fbsx7Amen6Ae4lIJY8y3+woGXAYXRLLJkypklEIiIt3h
U47JodPaIqoo236pQjneHZZ/oIz1VMfhHS462nyppuyFjVLENJYFs8NZ9TVWPcn8
vz7FHFOuu7hOFTjG5cV+Xwlftz0cSQwNdAszlRfAYUPo3QTG4si3SvXJjYzlAoGN
X12uXNOWzaAsFdODvNbPwtIvta22zFzBx41AY6wS1INWzyGfUd2vKXPiBtPWnE0j
+Ukx5SDjG0K0OXacfL43nEPrpF/dZ6c6L38Xl6koI1jhmb1Q4HYKbUxJx5btexIA
DKZeK2UjzH6KDeWx3oWeNJwFKByloq64KCAS6co7L4etCMs7Lxy3c1kyMVBfe+fH
qjXbs+GI0EfG4ZDCaSs+u+t/8zWQ5B/Z9U+kk6rSQo/FGuO159Q9U9WEOZLmRVZ3
5jnVq8B2FtEKJ+mk8wYpJhZSjkuPcNkuHFS75x6ehH3sB42ADNl/OBqnHi/NR6xb
LXglwyer47+ozwdmvxei91YvARyKafrp2dQMv7WL+S3lvjx0MEh+lE+26anskeO8
60Oit8C589gZda3Tv2gaSi3GzAiJPJw1ywGxxO80KAkih++PmeXEGiontoqp0xdT
J1GseSVNy3VSDppBAJurmmps7v3CGhds2xoLswF/cCB5DSMelkjrFF5KyHuOgkrV
siAX3oZxBxH+DyGq4ITnDueIuP/Ussz0H3/xCQZTElN6xBEKkNkiEE7D1F1z7tgB
0aGKEk5dLUc10c2svBWg8ftDUgoEFd4b9Gn46sElGIxrAJ8DR2BCnQAN+gmVkUTx
D69D20uLYw7wd15vt5PSxJaROwy2CSavz5Ic0KI08iu/Ml+DkyTWnDiipFwjHtpa
lDJ0i30xXQhG66jDtZ0GeWL7zE0dNJfSmezZRt+6GsAh5+6CGUm9epJCXOGGjrIT
g0CROgfYp3KwHp3LtTLtthveOA/fbXDBJF6LHg5xNZ1EXh5uGpF80sSYYIdAmigX
Ybf0yFMzqV+DimIRwrV4zPcGbm1Ec9QsRAOyaGEE2/QtACYc7qFDXxk7duuEBrSh
Awe8JfHSqeoh79IEzi4EI775nu76ZMP14Fkx1M7m7W7EmHLda/ePHITWohnnF1wf
rtV/0IWwEWgxUlav5Fc514213+CKOnXr0G8v/aIZXphHu4EkPwb71+91AxDcBo6Y
5BX8ar/o1lq2CrV4LZPz9FpteVnOzrJKHiGZ7pYOxg+FtUwQ2FRxCb4zxr/o+zKy
i1f9V66R4/YzvJgJvhhDVZROfDzcFysp8GhSJfVoXnK1XzchzmfPDeKeco4fLNrY
yDFGtDEMu/q2ZLR+8fHwe93CYxTElgjg4RJsbmtIepF6Jc+P8d/dHNDdbQAiZvYx
/xD4IWRzzBBxuuRsyP7vuyYcE33+LFgAn3w5uKgete0i5OVrBXMJDkOBlGxT4Hgo
vpS8iE3bGlawxxoTFe19h+Psh+oVaBfehjqoHPDtcU7qdxgpM9lGlIkKz94qC1oD
n6a8q3sNlYSeMckDUMHneuXI6QDUhpulojXYdaI0cbzaW0Ojozf6X3p35fY5s4TO
oM/wzY7Mf0ETn6OX/TaBSXtpyZpnOWemi6q6fEYQw/s2wZ1rmNLbrl1ur9ge9Qdz
NP58Nmd8lXogDHbCrV3IlrfmJRVP2VN+L/LwXufyaLgmfaPWF67/6NZese8tA8/R
xAvP7k3uJ6UC6+/v3VgSBjuQACcTptC3t7M2a+w3OWV4h8c4FiOZXJv+UGapRMAq
e2Z2bbbvR3coR+PMHHh4PCkwtcNdiWBj+uQVIrBGAFVVfEEXb5gjfkKFvoczwhxw
IEEg/63biX7DCLciFjibSTvoYEg71RvOdZ0woctW6zrGYUFjMeMJbQJXszlbETDK
9QcN5hjHKyviTvdODFfKaQJ/apZT4eJAszIXFdLH5Lq9SxJH3/PPpysDU+8q57fc
jzXIAM2cDHa1brTeFclCDdjQCMLS/QjaObseNB7n5o2TUT1v9y3Lsz8LwW85pJ1O
GjWRRBfG4a4yfdOz8zpREgmahmCpy2Jd7FgCGMkFj1/eEvgK13EcoKHgSlsADCT7
piRGW0S/5mSfXOH/hIfJ0QA8UEHVKXwhQ3KkWeoqL1TVfQVrAu/5rndCUkgI9iZ7
nJHwtwNlCJk0AoM+bBww7C9KGoCCeIVckOoAjpa78lvX+JxIWD//ZHiEAZnX/v1M
j+4VMbka77C5fmkAtBxk5jXy3D01EWAC3Zg/51eJgwt7yFcdDTJMcvPYP06Atx2a
G5kHiJYRhrSrSI9KSUOyA1+aIvMzdkOXJcFsSEUhEAgjSY5IQyK4BM+sgWd46TN7
USBTMFJGNQzuxIRjqQcd5ueWj7rqz46DWdoPuwjB9UwGgf/HfM5Kl4S/FjMq1K3b
mbvYpplQthCfAYvx6Yyzc9nsm+nsdhIUeXl5RAjmKsiz0WuNODYbOcQvv7F3+b1R
q2zHzLjwpNDEXBDYSJIJ6exgoDyGe9hQoqMe1lPsWyPQqhDXWcKJ1jDJMPRPJf0c
qbdMWJfdyRy7++O/miJyBssffTPTc2e9ZnGDiSWdnalBmhYpkvoswizceEfS09TY
lywF4Mq/Gs4rSZ3aKBRZvldHRUbK7V3FVDYJ8PtOkcAWIWFNfBNoxPz5ILIWP03s
6Zf7L7Dyn+g/72GW8HzoESdXiSmRBmSq5kLkx85TpSl3KHktW0FMIE7D/7tr0yQE
IhMs/lnWBD/nwcU+nSooZQSkT/p0YUNBMHvJYIvr44pLhM+63VvpUKqMfisCtYYp
Ys714JYNvTTSzDFIG1IXaS08NCCAG3wL+8s0Ifr/guJJchGhHpyU/YfKramgdBQw
DzubCAYVg1kt3TaALLvpQScgTc+VT1AT/iuLY7YDS0DXbsVGUuXzcVkjDK1vP670
2wtGTjvxcdQ/z2F42TSszJtCK20QgabXCdjmiAg1OVl1Si97Oku0BPL3fXOxQkMN
9WMX3M38dylTJtjZGNjB8Pr1FErwBfwMs+OuTfQuUEFnS09Y8/14w8AuUAe9fBA8
y6GLEO8heQTotjFl/ACp4amAbMt19lmMfAK46tD1MG/qKUMcDz2dQzzkz82+SYO4
OAmbkeS+T4HYy54gpN4ohiw8XAHqv2A0EdXtU0KjrD2zJO+i194E6m4BvYfqQQ0v
iLhvgTfhsRaVug/gCypRf8lBymKmkvTIaujhZyQEVREZVBIg1kvLVD9I6DpFd4vx
jbSWJnWSNDjj8IfsZBVTg6sBoWVrYgywPIz6LwUNn544WjrK3bPQVxypwJtAkl1z
jNSdd+IpsVrTVfwiFhK50qVSpGDnqou7cLAC+B6PxlvaJ0LC2tjMA2m6jkAVQK4B
4WbcOLu/kVx3cZTYQ0bZ/xM3TKAIGQRoRLUTIcygT36u49p1zMnkwg4vDYrpjo6g
oQxCzKfIEhAxms+QwE8qYcoqT+binQdov4FGo1UqRyc9SC3v4NjeHYPpUADISaYI
r6TpsG54/wn+pGbhuh4PU+Quobl8y0QwBGNQB3mAI5yzXjRVwQoe5NfM2hIhHobH
aixitfqCVhkviqVA+upc8gMuDRuHLNPYrwZjk4kl2TfDqQJD3Ho6NfVs1BLalfl0
i5cj4VuyPWyTh6vpX6zRKKqzHpxG7MhcgEiBcnsknt2IL14doaQuMdb50kZZa0O9
QQu+akvJF5UrEuP/BsC+1/8PNg3D2m8mhhLwFcSsshtsd62R/Qz/8ijcDAuTn9qI
hwPLT1UV46h6x33qFt3yjShMBeOmFPSVi9fASrqXvbdwOY+GDmC3Y18SpIOyLwWC
98xu9d7FILPEWmnKnvz77a8cTQN7AXOvL/UpTJXfqbWiP1JfgVNrVKoZoDKJc6GC
O+XYzXdn/lR/XOweXK/dtcqDurEIelwp+3jBar6CbvZ2u0pe0lNYou0kMOtam+vp
hcpyeoTN8N2fz0IMbYrp3DIDvvvjnJW4jtbC4V8EpiIrltoyOadBUreiKX1evfG8
SAsPdYMxD0J9M1iBBDPMWCcbKbk7Mln73z00VrPY5EcBzD8Xh/6/4MZcul+T21+e
8gMI3xFtF+u4e5Beik2zlelEiMU3Z+mAaELTwmPIGEQRnKoOqC+0TSmhL1nupkig
b+YZNV9MVsFsZ20VTxCgCFt6uSIATcT4Y8y1spfTic/wEhsce6hpWpxLAUQpNQEk
mnwTtjUR4oQ/Jg+zoG+78elI0ZCjiD8xmjNqZ3TDwdHGl5Z+IIbvlFbG7OwMV/Md
ZwgxQxBs5eehZxnwfFtrOAS8oYOcXMts0OGz+XRgu/PGHXCB71czTY2ClWEJHW1e
k7QR/U45H8MJVh4YpxzW9jv2ateg0fjwzA3X+wRt4Rxfub2eF0Y6C6w+EUTZN22v
8sDdNIHJnPqQJkcON1bAJrXeLgMYcLgbcMa8xbdW2izLnev93yPuVjUEw0fcJype
nPzfc8dRoy5PikYeAvylHK8VRGySlwjSEa2+8csJTBcH/SKcCvTwKtAIMoP8Lhr2
xnq3ZmYjUyveBL7Z1DmnLHrQQ5FbihUADtj8BIceiSJrzJDJz9lfMOXuKruqkOYL
d7F9Av8lOl7pOHN5+FIdNqkd2gSiPlNel7y3sE/uBdk3UqKPsn1jdZD1my5ZxnF4
vxyXZnjexZqriZXMbxi/9AoOClQ30li+yOOmw9unhnSNG8UvTMSo/7totpUv6N9c
HvVtUgy10LCJLBJOEZSz1sa9eFyYgXyM0Lkq7bJxcGLAlHqioZ+S7i80dEPJ9FnX
hOXEGoQk2iZSi7SWoISnlNEsUFufHZYN3FRMnkUCla0R9AO9GJ5CWsrVuYLQyoDg
Qc6APcA/EMh0S1ohfA1pcs9aMekB+0lt/wkpVenCAb8I7Yyb8TIE4LA/pJraRngM
eB7jtoJtSSNgfi4aOGBU6396aNLHzm1XU6STEp+OrU2Uo6ODzqhonjSu1yYj3PZ8
/+XXFijG6GrkOuqKw9zmWd9dx4Zk3uVl20VTd7O9DU7OuIOLaL7eg3cFUKwqZDYp
XubepuKdqu6WWuPktBXSfTbMVaunbgWC8wAo302+GRYKRH5HnouwJftq56NyLIQd
+mpyQQloA7uBp8ivTv0PWXXFf7qTeQk5CfLn00xhAu/ijS0ZxUrCwMcV62aiKHpv
T0gjRAL9DizEN1AkqWCyer4AHQcgshFfivYFSjFHInGH62wyg4w5sQ/mh9WJk8q8
X8T17rUkYDxIFGPEzvcqf/g320YHMT/sBn8lIh+mNWlesd6djxtchqsz3/Q/iNM4
`pragma protect end_protected
