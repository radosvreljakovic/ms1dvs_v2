// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j7ZaYyCHRJzObR/T+0d/ddzdecIpPHZCFgRS6hcfXnLsY2Uj7HwYcJ2wc7Kv7vL5
E60kSzDGwQ+K+PxHpXR1jzIJphmf73UoNUFnqfX0inZdKoT4HLkg8dYIDxng8TS/
2sIRGAKHxR8RL4uxHklxVu03mhHN2dXUVuUFFgj7ZX4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28496)
e4luY7wGJVkt8GNj2Unb3c8Gzj93lU2fIUZIeT9YQTTDK/oXLTKOQdcUAv5SUYz3
PwWoRmhIoQu+ED6itgfxzz6HLhYRb3gaCGdBCwfijHKK8yJpCCV6l2yAY3HKm8RY
SyF5Q5kkFI5kF9/Kjg3kEZD9lhzSPZQxwrmXwNSqs4n4VcYF5jzj+jzbLM9jtGtQ
RTcEzwqxrrred3MfYoTJ9q0NCxzO5Gm0s9G1Ixq78od38TY1/xC6tdRKOIvEp3QP
Miq2t1WZOkt9Pm/KzxbAVULKh73zrPQZiAOKxHC61IrY7Mu0xZFkaz73eZSv3YNx
48NaZDrerTmo7S/mhG/Sf1mIR5jnhMKt0AJzQut0KDYp5zo7vw97MPUPnVeCK1Ij
b4yOFSucypG0fsZAbKjVL4gECzhlpUG7G/gNvLo/XrP+Rlz0/c/4z8gGru5uyi1i
yXSARa4omMofFNKfJ16Bb61eCoeTfGP5Qe86IDSWJINnkg8l+sY/+MHu5WiwAKJx
wG0OqVhia/U+w885Z9BC4BQrSBsSL1t1J0ZSmrDhq5ixW3Gr+rKiVs6uxgExoqyY
0Bj9HhhZeL9zeKeSCCzsKaFsBIkDCrIxEfzZSA3mRNMd9e/W1gw7A50D/K8sPrQl
fg2Kll7h/LJluPyqfhHJqjNpg2jphD6VNWJ0yZYbHBBhWmmkgvA3Zc7Sr7CHb2Xp
uFdXCilUxeLFaJaTBuLCj0cpkusbnWcD635kDyTlkTJfy+qBmU/cCz9zATbvwezS
mJA1I7k3c2V0fTh7jZ5ZVC6SyxHbNSyCRiW+um8M32Z0ylp2XOGr2NRFpZvJKAov
0XnYH1Z9k29kh8elMrCRUVr7dxvsJq3ADipIIlttNOfVWp41odH1grjewOWWmpFv
rzp7YNqBd0whLF/fTmWxDWki3fsyd3UI0o5lGNCmipZKoulQrsOnHSXUS8cxR8dx
oLnGjsvFqZkPEmQZ7VKNczJ9xF05NhGIUn/bmpqayooT4QdLl1948cl+DP5vr6ZC
zKvWwxLwCjJtaUl+P2kW/68f2sXLvHG4BB5AVDOwgcv12ebqAS5f7LkE6XeEMSL/
eadVZJ0DAsy6E1iXT70OSjWVj1mIMc3D9fIJhhLttlIip8AiBwVkhlbRIkascxzn
UPXTLP5y3HDBwxuuPccWtRkkk4Mzjx17wlFpswHVwAa0jTPAu/8zWWwBelxHqUjV
VwhB6MupERHrstbdM+o/DEjnF9vY/tugIXwCvzHuQG0m2amIItoy/jHWFijbdnuP
ixyzpYJq1t3U3lNOzJ7QAu7PEyaV56PbQsCXH74CrTJiKed8EN1whR1KugD1wHfO
5zrg3TclW4WCdxfR9ltks4JzBu1dyDRUG7WWcYrVVMErSd4hwGq95iJj9NBgiawi
zpqByPf3IyFu6lMIcZKACRL+ufJm0Nge5vXfRqlD1wPl2+sPxgJoB0C5VJaKvcqm
9e9A2V08jPZbF13uHAuc3SNTnjem8hirqbgMqcEo3lQlWCoxKOW+/Y9rMJQMiw9E
+Si057xl0lUVsKRZDEuASB8NE2hzaQyk0gyIjXqYt/3n7Da9S8DbtoyipnkRmrGT
8cHzShv496nG1LcCAjV+z6fiQZtKIwZ5D0VoOXzM56m1rkRY55ODUmooYwc/3MEY
5Id37sOTcbQJFC7Nq5DNGIp0BLf9hH2ne6Nb+fiy9Po00VgmdspupvxU8N8ZV7aA
Q7cDODqZz8v1wUP5DEuB6wpm5v1c35mxdCwHNpqJ7adb9pjm/GbgNCaOFiLb3Dkr
VAtPuSjEHsFLZc0j4871u+K9Bt+7cQPuTm66KZODG2eP2pFAJULr9Fl4q4VOzq0f
DXoYJKv8a5PL1Q/bCUIjqkeQ5FzamVSypOUystjWcHj7h+r7jAehwshyq84xOIFf
SCPeXU0xPvJMmLcQEP6f6cMm+sLWf/uhsoLY0Tra2kRQN97SdA1ERTE2BOfcue3w
T9MnnMq7b8sjEDjr4keSL9584OjfFukp/wSw/adkJAcfJlbIbd1ZzYTPrpavC9iQ
M3vmFO27N48T524HLlH1BX6SajEh+iskBZI9d7N8Zsrc5x0k9kviXmqb8LL+QAUf
KTd7RBQ+mLdredTXMgYZcR6LUw7bKp1p0h5EJ0TdWQdStAorP9k9X0KtI/+vZNbP
LpZ2To/ljfHl2wBjUfIuOeQqNrfWKXJQcIXdXQpSUPGYlnEPqm4FgRtIvPxEFQ0y
w/ZolLNYGRRabRq0sF3aOgscFKu3jkD2zAkJShT0DSiMdNI2pDgkS8W3vdGaeAZZ
xCFzeDpOoev1CFBn0F2LdYIKsR9GNo5Vhsi48NaeSWuAhH10E1zG90W27SNYKhyV
n7pfyXMjk85tsJd8ZFSC6pBi7X86L704SQYVLsZMF0Y+hIHOcXBgD849P6DYGmKb
VdPvDzYwFqklQc6BGOlKMBeJORYrGrYIOlFwtGwuK3XGPeU1EjGamHGdMePAv3b1
Csnl8N0WN4AtsbtC71zlWZV2n9EAvKQx6bt69Isakw7mE4kz/HBNqBh5H92epmUd
nEXjuvb5t5OBpyqrH+ZEhZ9goYtbPPgVYB6gFXp+7AZ768pSHOSD/6LwVDp++/Ce
75l28YI441ZUVYp72S2Dhy+sPqhMdjBIHDrJRJWIOh/Y8Rmx+hpbc7CwYwR+8eIs
2Dln1Udy1DKkGnl8q1NOuZHouWZIB96iNZNbxfKzkVpQXIB4cHXtFlwmNQHjUbMF
hO73zTvegSAa+9qJc1ya/9QkW57HRZjcfjunuDzumKHZhqtTUPr6K+960Y4AdjB6
2SpFAWY0+L2a8IYedpFjXnl9KdT1WI6rWaWje/n5fZhDvqqynjQCTPfockllWkZc
PGggvZ1Bnpcs8wdEhg2agavrFdomG9yag+J4BEfxgCUGrFK24LYaGugY0J77BFtx
QyhVvsk01XPGHHJLXU3PY/j/9NqfNNo11E3zUR8x9iXmH4rtCTfGCOKExUpzYgdp
c+bMdhyBZLeWJHPY/we5S+I8/qs/pVEPpj/ITPz6K4juSwHdZq0AFW0T16AdShYt
gtA3on4bEhFUre8n6iAHAM2L5ZQF7UKH93wHCtJgIH1Yg8hMQz7Z4S9Zq5ufAOfR
ZwA/c2JpW9Y8KWn5jOFJnP9yJH9kqgPJ5Ll2dGhhi2OYnamWDjAlpUCHjs0Up/T5
4TYr/ClFwvm4wOhUdfWCCXqmaCdCufi4jlQUZ6CyvnCtS5AcQhAZgczWnDHZRcVu
ty+IFzlCgyadynWk8yI+g+dgtLTihz2slq3VmqAaiacf0PwUxKGeBfPz7idMrPCb
BHDg5axhoKO2qEkO+tn++5CP0tMLzrUwoH/a56/Y62K6WYOsL5IOsRY9wZrhar2X
rs8e5AvJTSaRGSIoNb77yt9FmUP4Z+Er92raObU3+8EYnmEJUlurCGdiQ/2t2l7u
wMrBPRKLXaEwQsnc3oHPIOaNfbIeX7ToTNGqBW3N21Jnr487bb4FFdbGvV1J+24A
BpvpJsJi/DlEAUoKZi/PFhLLYe1jYQdm9UjVjX1ZwYPATsFEeLZSFJKUgrI1FbJH
BoIsrXizLipCZC/Ol4wrPoOgEjdcF8DJ/l0Yt0rPUKmPFZMGmd0t+MayHmAhPd1c
ce4DUWStwaAFv1QRjyoBMzdEK64HXtTKckk6JicB3bc8RP9HXlS75HlHBj6g4myG
cgJtUDb7aL7OrwZ0++q3kM7m4W3N8UcmqcAioSVv+sgpSuFYHyhjtQobscH3AR6u
sOeeR5F8sziM6e6AyprYSMkbhikxwSSZFqd+4FHtKRrzoJ+aPsyDebDmXCofkD/G
mUH96SiUA2sFS4IChd3sgVH1d627YuwUHi0elV3HEI9nh1uiJsLga+U7rl7UJv8W
0rBwb/aNlWCXVIqPTW0b9IQvI4pmJ4pxDRViaKu5sSgDiqjqL07fV0A/O8QVQI+E
tMDwy8xMV0Pfvk2LV7cdV35MJ5070SkJ2v2FJMFgojJtHM2umrFv+x9p8oY2MJ5t
Oo+gkrbKIx06hDcHjfCtailYHz3C5WLc5rLp1D8DhKuBhWSTraYRteMZRGjdV498
06GMxzk9ICQbnpSxuguyH3/2o9Sk43vGpxYqjZwcSIpGoUt0h4pfuAi21zbg+teo
x7mCG7slHX8/pgllYJa1bEGJuhortorLSomuuArkP1CRtpF9N5ya1Ui/rudsuAAZ
iB3XOm7/gGzNOW+yBv8LUDL5rxqBHewjs4CgTvTjVapIaLLNYC7ImFF+Mlm9r1Sd
1/OCVHQDugj76sWEL0o2ryC+1jvhcmLCqbTjCeyMwVw9y3RIBsU17S5ldUVsrIfu
3iUO0x70SOj1BROVweGK1dkEymwmDhukR4GBhF+hJYw1VMmxNrpsnijJQFW/77gn
v0TsfOnKcWvYyJ1WloHRRUxthyLdVaKtzrL3RMpNbptHCco1l877oiF9qcuVOhFW
psEEBHNc1Zc1/LRQbuk6ES18Fb+cgJIQJkERXcYxHdL8haNbcK9rPyNrDDE/iY6q
ypCfhzaS46jKvClr704f6A6cj1lAtwV5Y8OZq8B9rE+k3lsd5Zewh4Vn2rDI+Hgi
XSvOreF094nQmg1ZJm7CfZN1m4/aY2MiwL4LjRtZGTLNRkRHwW/J8K80W4htB5sD
cgbFmt5fPnu9wERvZrJH4cLfHydOJS48TdwcVTPj2p+LJqLhRAzk5U/w2/FexKnd
DG2aY17hyGf+ocZk7XTszoov36TD5iXvyqat7t6aaHYIprZHaq5FYArQkntgsQlH
RTFUMqOgLj0AJDu7KnalaqY3Fbfm/8eio42JBoh+olSa3CQJw+/9j/IxW9y/0ICp
VES+e4s1J8Sl0fGkMZ1DG5Liv2XCpcfKbps0FFtTBlxFCD8GtsCa8xH9BMx+paOm
fR5+Qc++cA84ZrMXxeQeNDcUIKlu+l1907rpp9DDHZS6JQyB8IH+JCc3D3VH1SX5
xoC8PZCNP/TIVC3qki+q/WF/tUMkZfD/9VOrkuxYDRYNsQdVqyniZUaKGftXCJ8S
udNMts2LyUF5dvqaKvmH119wklRXeOajG3P9uyx2GIq5377xCM+eBPjSFg8ey3xz
A1Q7+9CGWYyfO7Z6GzBci/PPrFQ8heCzNw1oRWtUKwyWQXJh38Vw8FXRX8iVjd7+
7se38nurMsXS7CpKl+xqoEsFIG+16NnZ0RT80592csIJVRQf+8uiiNxRvOxWZ7xw
WODsRbKPkqAw2XUWv7NGBWu3J6Sr6ub+oCnUy8zT9ijWmAKY7mkMKYy+gnmukBdI
lleC6PZex2qb+3ZhL71XpgY7cy5Bj/D7dFhu9xjOU0pG3UqxzBZUECnrUiK56BU2
sridJ2r8Wsf1DDCi81AEnEEUILrC0GlgauY/N6PWW6vZUdFFzUeSKaD426CKvf6x
xma7/QDHJ+hnfujC3Rlh6nvm637sVUjDPSXtBjIP0djYv5o3ENt7LcgyXydpTh9g
oJ2SjRLGeCVwkL+kyha1qht8835JK3ktj344jMO60hupwQbTYscyJ4fbggtwJlAp
jYFOO9RwTEjR0B9XK9Bx4/ZetFOgnR0L9YSvDS5ByXHMHrQy6Q5g234ekUvSxt0b
m38Q/xmIAeQ0Sb60wJQ/GxXnJp/faCev5VpjsdNfI8SmB46PoSuvWiLosSGAQked
0fhafSL+Mjvhk15BmFQm8gK6AC+AZrBk4dMpCciKrVA59K8ktnaRZs9ArJEpmLxz
0qVtscNubIRVeh0uczoIut4xydn1o34NT29/O2WN8ndlJ3vbTjsth16DXmGjISVR
iEeBTKGhQR+kwbvtP0PPLSv4svMFxHC30u5sHp6QIpj/GlOPvpi0ylx5n57ADZQk
fzF8GZDM2LPCYgfOjQJd564OxlaabTBVsWnux3NIb1OaXtkn0WFdKNNKdv/WUupq
9TZBragM8Kish+gR/uaX6p1cLdjvvh0E2VIwsuM2EbUvsT4ByIfw945Sa9pYmL5V
xox5A/BrgJBMAtVqtjxgsPHnBtNHCBsFpKQaUhUvT9S649/LqmLbD2nuE6WFacnu
1Y88aGCLVlSXYHzDC/wMrGRS0UFXkyiD7F/49o9QG0XA5g6OEdE9dtHm4ZzZQj6U
Md8UyOv/kGwJ9LVVv130prA7tg6O01pFEWwBDAfcljDb+ZwFox/j57iTYc4adC2d
wskHCjg+YbeZkhEK63sMsSbTFmLsx1pS0VpxCZppTAaO9IbND9R+Pb6NegFmIlL2
tbr+Ho04IQP8Bl2Fk2fHv5nvLaeVSYwZuBWXamS1mAN/IW0/VQfshu0rxDd/XNhR
i3s2aWmBkKTW5DzOqiK5t4fhO/1OYuToHUiVhWy3rBfZmkoDxSHziJPS4xm7u0+V
3WbEt627X1Nz2X64PkJjaC4Ae1TwV/Q9aQ7/IcaYPyXustrVr3oReRlk6B40ZQvQ
n8K5xZxBwIWg5d8cm0L1GuxoRE3TtRKhZV4pcJkEQwK/oq+bAi7bgDYhrKVBO+AF
cNArZ0YpstlZXsAfzPM/CNys/IJP9Tt9OV8CQzO60HMleTC15HzKLvVGq0ONBAiU
w+1pEEucZ5j6r1YT4VtXMkwzoVp2TzNb+ka+I6trBa0Q20aScg4AMxiDE1B3J/Il
WCUuMcrzBa6mG1nmz2yHOrgnXjbFDiMzDmwmEFq3BJfDFeEIra5MB3DPAY/VcdO6
xd2MRgWLGLMO3BkOWWr7uorDidpXQ8issCP9Egg7HoH/10bcEJmSh4MQ2FqLRCZf
wuCoQHC3hgXnRqkNwmn79tvlt/KR59H4UiaCeoAq+ELmvhIMtYdMLZVtIaFzR22D
pZU/AZp0uHoVI8dvv1/Vk0jei55wNMEI73I2CMW22jIAGEpeO8jAU8FfqohvWQEJ
7vn9Atybzu2sy3q7+d+qUu6aPfFSzZ2uK6wGJzF8acsJvp3MRuqj4zut80qjZrNB
U9ONivkIZ81oUqZrGzFpZUBX7cfhink2+JBpwVSJdmoSumIfwZ4b59dYjUucgCUK
O2bwDQUVUT6O98vP5RyOqiWfvBLI93jeePlLxqjTCjrcSmBn94DnvcerGrujByHj
BMfsje19FDagSp8g2Rd0GMwGyLzcmfcDE5Chfcy+MMilOJfL1pgxeos2Ly0isOnw
xJDCg6eSUrrn1ZnR02JZQ6lnlK/+Z3FLsj9pjalouQDQLsOhcgZy+YRifmG6Tbn0
MfOtBRMFue0CCyHAyq9uxpc3PFLuTM2DT2qNYsKd4b3y4t4dLZHwitEZTiPhi/lf
f/nYbhudSNhk/Xnr9bxI+5N/64UgTg2gejx3eL1Ci/0+NWet/Ef+bmycTtjU1/YD
hTrjBp62YCIAA66zLnO6feIptq49tfoKqXEvO5sgjEYkuprXOHsB8NJ+EO9Q7Lrd
4EKbhVO7/f65y+J5NlXtk09JJf7YCvRuS4H1rsz84TbozXZ/v1Xud0Hz3na6zP+J
rFIYy+VPgUVfTMT+LS4e2zuuqNuq3hWFSASCQJ1HMwbOIP+6FARKICvrRdn0q+2e
xRFMlmHutXQEXQSrlasZUTzHrMl2/sKiod0nMOF92G/QFTb8Ic0Jrecy3JVoKZ4H
/hUVVaUdypJTZidkKBIa4mNV+5LFEgIve4e5Xi30MWwv+oZ+MjOSUKsanVg0OBQG
rg/W+nrYH1iNBXNHHzfIaO7jpx4Va6eVtfDFLctH+d9U4QPlgFINOfAniCz2cYaY
7/phYeJVomsuDK61Fc9GbmTFjQh36oqWx4mNv05IDP1a7ZtLpat1ZnvOegMYUWf9
xl8fpyGkBwRKkenVpuJWOVpbxdsrBIfkNGbXSInWMI6Ci0VVH558h7EI81IewM6E
7gx+fU4VMlXWo967tPFIjTVSoRyQqcIzXa0VLGSVTEGIjECk1+sRw2OoYlybOWP8
zWcVOYQ7FW3mh6szyOHISv1y3Qu+jk2b+MgU7WBICjkhkgThFcDQx00FKKMojWIf
2WbE9VR7JrTj9IuoWMaQ6vSPyWUgMFtWMv/RwdLW3/1cOd++VCPoGx/Cxeu4/Nd7
xdCXMiNTUDYFZThEhSNoFDhT/TSbDHlvD3z14LU3Mnaizbc3X7vxfoTTt985bPnF
IMREU1n5Slr4s8NNE44QwNT6Cc2FDm3ypaj1OHk+PFH9WS47BaLZjWDpn+oOJZYD
2WuwpoV81Xz3OgsFtWzRuJPiaqczQuAm2JZgBfa3/foA4ZabBDRFsfVUFJmfqpbW
RzXX2nQ1/kDmyFzV+01UcCFBSrFwxv6NG1mphyeaxiVS3UDuNqMPFPIgB8LFYlZH
ta2LO3ENunqbxS/GMD0+DyZOUV++ppErgPBZEXnG9z/uOCFjKtS9w67fckyIrTn8
ltHtDDFwhEQSdwn7evHnUhs0MYPIniahLB5jXvOZG47Cn8P4nsY42xiQ78MKXN0a
rpstIwiK51JD7wAJ+K7l3ELDaOtP3Qg2fRNxvhSR63iaSsgeLkUxDSIYkCeOSUMd
iY2jc/EMrLzZ9ca9PfNNMrA+UDwAWkC3WUDLp5VONGFxZTJ0xepeep6NgFstS5Sm
rg6C3vfnaacDjjBl79pcxsS4rz2wX6FQTzrImgBFjEPQvWtt8Mue+55gCTarhDc7
C37kQdS6Qm0tzx52XitPwbsheIdmJtsTUDn3vkzfuHvEhN41yU0twQrJI/OgJC2t
0crHDomENlZ52xYhNp1yRU8Cd56f2sK5pTxnh125sBLWvGcYyEhW9EAQV8cZYDGj
PF9p0AaIt1g6kjrKzIAzapwqlafRM68PnxlVPUT5HpU18hjkhcLLXvY24mkR3ah9
P5OkMg0tE6rA8aghERDEPlI1H6bAjNeu1yICibZ2EcqiWa7o1N7n3917kIkHJNcl
Dn89WXqbL6r3y1jwpKPFQGIs6tKsPpqfD+JCGmTTbGRrg0yQ1cGRtmA3Tz6OGKSb
Drk+fgLdy8LtAuWVxnd5Uk3kkdZQkEUFaUs6uKeYVwXeKOv0vfUiSGnSaOx3SG5S
Oo6ngqL6oBNkeOwWTHqLoVu26BZPdHMTWoTdjl86l1T0G6T/Zwk0Bgba4k65UMue
62zOxIo2HQlvAbORCX88SI+91CFe6qMIblGnJwUy54tBEqBXn1j50wT0WdeIl5u3
nKJh1vgntqOJbmFTUKFTJ4FclkmFH8XnWEFocNQGR75GtxQ6vJ8vxqy19t5glU2+
YzQmLf8fNKtCOt4XHiblhKI3ItwRzSFYSpj6J/zViJEy7XhBcEI/XHg5c75F0iLH
fjDiFKAL6GA4ep+EXA62b/g6Hbx1gAvoXD6D+MGZ/knVBiDCRf0zhieQbk4pPUK/
X3jHqGL31lKb8NcdYvDjKJHJrFeG6Ko2L6yQwxI79fT4efXq+avfaCZ5ik8erfXl
VuJ/66D1321RVSjYZMVXHUoLk7xHhXULIvfrrhn3ehBQWG0hAhv4/bsaHIdh7EKS
y6u9IEPjBd5H2VkI19PPqTD68o7sKAwyw6791OnMyIB3fzc9phshA4S3Exw4raGp
ZyMZvwfyFPsiO0dtfzoiI5GFFrRMFAJG70U0RRYknOAHkRt0RTj09HwNPgZUKTcc
kxKLjxn4PBuujqK/nh5BjUmnOXpz3sXQY6W2pmHrBlQ1vCKeBJAcl3yoGRBhYixK
jxVG322Rnb7BG3fiWoGHLr8D08MEPspvDKRdyVOlNZvhMcfbfneogtO2heHV1lqb
1DzMJfOn8Zw9mFJ7nrNs3eh4ICUvEsRf0HKi8XGXcjNeHGwBSTyjCCpnwfg7bAct
voW4MfbYpdXNK0U+1lJi7xp8d+ssDyD3D98Kiqs9xjeiD7scZ7j7xw5M3pc34z07
MTKGiqYwZzGMNmMNr6ofSztu72UHpymYRlEyjxFDwcrph/txYzfynlXHeryeh5oP
t5adRHrGRFOQZC7j8JrR3A1uO+VPsNgFPLJRkDHuhj9whARWbv/KGxoVmw039C27
yroaABeDxpHdMLgTPzb9VMNF4zqLWJIg6i5Sp0EYV1Hxvr1WniF0UibQ4U9Aq3xC
MRh4YtqQGFkacNt60sXdi9UUummUOV9a7i50N6+3/4J4kiYSGqsV8Zpnssc+rkao
PFBbz5g8PHyoicbXh+6iHZfmALNF8+c8OfMMZCwk9/NgRG+40Dbos6o0wf0VdJcX
UAMm5pjR0UlhoBGDrVc2UFuaaIIHpkcZ6MbyrezVZIjxhmFXZkMR6LzpFBYU1L2b
wurGWElb7xRyAC8vG1y2n9a/v+S6W0/L0wnW6saqyZrprC7j+oIDLlDWDcyv7XsH
+5t9gWitMNht884UuSCLkyshYJWi0pqUpRTuKpHHYjksScmeTQ5S6LxzVbTqU2oz
sekSI2mBRQBf/0fT4+54xWeMVT/1fBsmULBwWJOVIhDHPx81j9MzGa5jDXTS7nq/
errtrELwMrK8zRkyiZfxCF5DGR28doVjX4WM6pNDgseF5hTNkBy1zVHv8YcT+0mw
2j29MTTQmTRW1439qvZ17haSMnQPG8igAMbThUwTjvV56mEPE8p3cCHy5wdhV5RB
JvdTkbA+O9fZIe3IQj5eKuMn/kGiUxQGncBM9GA2Y+vvzLlHTnszkZDQLLVzrmw/
kB/NTjGX6AOQwDY6KFhnMqlZ97pO9mt4tGXe24X2ZdsHNfre/xMyfacROyVQr86t
iVWt1t++sWU6pg39nNMzJ2mh9+qkCIBaQkKwqcrw1Z2cVBGfBw/DH8jI2Mf4zs2d
dwp4GtSLitV/2+zaycQ0nkE/Gs/JwpdiZGshWykRziZ0YvH1oakZeyFitZFDDdLl
JFt2bVpQubXmX/C37CqYLPs+jnOKm+LNZFHw1ck7jogs/WH38A6gBbKBpVVbE8a3
D0MSLDvw4j5qS/D2fzJ9bYDbJFI2ndyVGlQE6d+jfLP9C98/p++YWqm1Xn8toYvw
qTedn6Wt8ldoChLV5io3XjgZ5+MoacAjPvKk2Vd7dKLeKEx//NDHct/SRSmoYKDG
ed/ZCBV8PyMF5wwEP64E34KyL+j1Nmb0RsnFeD9rR7QBQyU2Mjw151q4r2RzmkUb
NP6vemJ239zhPQNwfW65AGcfQBwvnw6FRnqD61j68T0HETHwcMjXGssXowkzCDhW
g0YoXiKpiy6Mj9XcmZ7mAxyNUs94rKkGv6v+km13oRCxswgFdmaxScZxszpnRosZ
y7efHEmtEmUTrn42ePh0nFjiwNAjsAjGYozEXsVjhWs6spbBkvX58u0Y8DFuN3Fy
tXhDrFrv0yAvHqkHCyQfGe/Wyl5I7drXmVOEkk4a4EbqJ1LB/c2LwYJ7Q3M/5Djz
8swiedhYSYnsWjQOHMAALWbHpK74BIfllaH/pAlgWzHAFKSn1wk3sNYzEUmkh2xG
1D/G3EsaN/dOj6pU6Ife24t+ojUviydv617Zskae9nzwkDMvGJhl/nXJCCj9YMPp
yrPuznmLmRP52GCPb/Q+i3ktHdMqKU2LG4birvHUD87TB3IVQ9w6yDBHbqpIR+5j
gM1TWo4Jtd9hLquVf0UyTq7o9PBfeT/eVHccM3I3zk8npdAlOD3gToICKOi6/V2k
6HYqVeK+EduwKiO13S4zFcQ1kr9IMmbxMuRNC5SmUZw/N9OZX+O6hRuwI80m+85s
9Z4Ji3egoKiSQR3r+s88yzhg3NoQ1WOSnAE3Lf7yPAKP0PA7gg/hmacMrn2eUrFe
062wqsnTHuuuyhaUxQg+tITx/eVNbvdBG2af374PCxakZ7ZVFt+5d6uf3HlEA+T3
49yuPJLbyGsrXKI3RawOzdITMb4M5UUF9o7loCwICvwRY30FM+NsFME57QgSox2+
ZDNWO8BwgTkLbOFXansE5az1YKkGCFvH701kmodmnXehHvVk+d/nmeeqDzHxZARf
1J6Jsq8RDy038ebG2K7OlGkiACwU1FXxgygv4o1FvWIXACaNOB0zub0HVr/vLc7+
EQ/ojTIMLkyARG+jo+2q/fdkXtgzf+99zFS+NQ2EKnXOIpY3Eg4LMLOQK0Obw5Um
V62nzAw1mEwDSnO4oS7u8YwnqAN8FGO1DQEHVupVSLFw42kTMJHhIW7o4//GV5sC
0+tiyCS9owjzQYvDoeKOF09WJUmF1TX4HBQW7k2mCC1LcgUNpdFjyUayYMPvkHxX
s+VOIdkblmuwpRTZWQJEU9ReJAmrh9TPqtTHcMRjWo2V3XQwzcVcI+rkdAscJWgh
00Av+De57tXpUF8D9b49k/48gW/+WQIo2mZ1K8T5tdlKrDHSHi6T88MpqmqR5CEP
F1hRLYT+pDWLHT5Q1dfxl2PVjFYpGjIfirkRDudkmEUqNnZ6ylFQoMpkTMTBXvKS
dVqrvtDdVQkG9I1Gwy1rzrGZtSRlEEM9OoE5QfIZA4MUN8Gb0CiY7o3/nqCHtkj1
+9oxxvtaxIqSp2v9lMe4CFRSyMS76VHca5RFehcdyBfWC9qFjYXT4aShPpE/dFgC
poKNIjHGyDF+ApgqvlHJYuY5xxfAIjCdJ7SLJuGb3/QHpVocMVhkLoyYe2Ppj5r2
rPnG3cLG8wPW3WypevTOhrOMJyiLc/GhWdbCDe53OH7gVkYeK8bo2Hi7q/7SvnP0
5wCbkdPoM+QfXM9etSanLU9JoaFnip4kKYFkTy7fu5wljTOXq/0c+I1KMFDEe8Ts
63x6pFsIYsEzf8kobwJFSTuiFQPJiLVs+2gakU7sfitsVIa/0PGpse/ucl3ghTz9
nqrZqc/bfvAm6+Ng1B68iDA8EqRldExnOB2U6dTaFR+p/uqdxhHcg5ro9zKLjIYa
B4JfU7DZnoHQG2VAUlcuyBdWdClGOmzQHrMPq+P4/wglXlpyMVG3lJKqKE4tavmc
pykw198whCUYOAFiYiF1o94xt+IfTiD8iTGlwSlbNYOJSj/tsqHTQkjN0b5I26UV
AO38YbCA7I3x16aG7XHDQBZQhhaZh9eGcSwFMKKrM7t13qHGJ1Yux0NjQH5Fh+0V
ItFb8DbmQLnat6Hy9fIMQckJxuN1U2euBJtIAjdYNTEQ11FKS29cWDRUv4RfjWtY
1K6c1r4r1GkBkH05FHMnwby7xWQf3+8KUCmjT6vNJFJAMQ3FXEa5ReT1W7XJlEb9
znYzY9cKGF9LNr2EZIYq4ANJ4UKl8uQQuMAlXQgSvc/mHXWZikOl5YMM5C1KDe/R
C3npq/8LbsEUxw6463mWCvBqiGKgP3HliS/SbYKfxt06OucoABOpcerU9kDuOPQx
4FUgkDNV7kkuOFC6cOIsyafiZeJ8t4YemBhkgDQRMdMw0GY33l5NwcLD2WtGMooe
z8aUl+kGAqoRIWtkCTfqfBXcUydBS0Ot5MTS1zMCOpNPGVrY+FRwKXoPZBaLzCzJ
4jlALp/+EdxJLPVOntT3hlk3YWiZu718JVGfzPAWKGQMB4NMXGF9jpCq60RfC4uf
9H18yCkfeq3lKoHsnja0+J3cCF2xKOqumEaM+YUTIhcq22FEPR94jmxbq3+y2CZ/
LBxyU9d28N9OBso31wgBDbj8u2z0Nc55vBtypSBxVwI4Z4k6U5HAKii0Gam6HfLY
P/sSllTLSNm4o/WQnlkHx8D3XgR7RWScKqf1IRS5YbV4axUtF4jQ5CVf0TVMz/vv
1n7Ie4AqDLXjFT/UzRQ/VUfJLXElf0DkIcC+1Gv9NwQBvULazfIxLJ/sghZe3NZx
HFeJot3Ca9YsqpjyLT2OffQunEjzZs5UbdjUhjo6pjhPSFl50CCM+218khKWHi7s
3TkAI8zj8QsRkw6WqxXaICvfRB3ICAwHF89KM/SUkESZHZ0OcOoLX/W3L6j++yVe
F6g74zgv9f4dkTP3C/65QMMKp+m4wm3uxmI6JKqvIfNEP+gWqj05hzkqQUEyayln
EQ1Aj62yy9fUvzY5ikDNJHu+9/ZASarx+cqxt3OJR8WU7erIby6bOQkzQ1q6eQYw
jZcm64R1c4oAjl77uSN0gwVpJ6bTeqUDz5w93vWxSgnXbpXJSWL6YZVILLzPdbwI
w1X17dBADKLkKfysvdnY3M4ea79I2yea1e8vgAk1rTnyKUvgNRHHr6bDIGj9BtST
eh4DVZIczeWCpKU9/tA6uzD8W4K8gwS8o53n7o0M3lmvoKbbIbdFhRuHhkNxUGh0
HrNl4FO+9rBzbSgK90SBWaeVmOZHlP2FvmEsYhZbTAn2IGrZtOSV4oS7T6UGHc/w
FxtjhOiYJFpHgXj0MdsWVnWnNZt9uBm6b6FjK3zxkjbOkV3HvVj1ifC86snT3nUU
1w7HNqAR+aClYlEqAoodur/Dc4gauZWqgkBfI4oflY5KwKrSERhxV5PuE2rRekXU
LF36PDFE9zIV4vmoRZFVI/UuqFbmpD4mcIjWol4yqPNijEwSHuR+dNHjBrEEZzV8
vgt/p2shTpAAl1DOYqIUoSPqWWWVNsW/sPje5Wshdvq+RVv7f5qusKO2MLMdoASf
9Lsa2WrBQYjcaps/b5mgdBtcXNCpAWuwyzuPX2srZwZN5BMzAV6jR64GW2ZxCvkI
+l+vWiWV/FFKqKwlw0T/xQectlGRBIM66o2jazn41LtXc7uLqg1ZG97J0uRSQXdm
iA70Et78HL4ltpbbhb38lvf3+4nia3oNYZzb2Bdd3LZeTCeGAIqpnUA/MMMKEexk
GLXLVxL+vqxkqZPH2qqRostOQbCNm8We78y7KRPGzat5BmWWFFCXc7cIttdmBWtP
1ud2IZWKqHNwfgOsjlZs6fHNRafnCTfM0yMcZBrBrcAz3sYqEhWZzsgBZPJUT/GN
F+V3A0/QZtfVeifS7RIiBLN/uA9h7PY/1+JbWw/UY6Ck4VPu9/70u6LSMLimriq+
1FRwcjHL+GIdknbomANXm1psWodFxr5d2LORGQZuMupp2RePTKLIvNE2kjTlFacG
HWfas2+bCJ34dYaGJGMVqvqbxbVV8HsnmStNlLWHDvjJMp2jf5IvveHM5tU3ji9i
tPr+Qm/Sce2QBTIjNdHln4ygHQ1p61dKGJcYlMvII0cba30WEb5x50gk6bVXiXI4
eI/0edk6Zn11EbPgkv7PskIg8/W3imLcXz0g1BBxpiKNfz0ovhxynADUrIcFwDwT
crM2/mKhvsNkukKnHHsdjKIr2VL5meOrX3jDU5DsIhqqeKinOQ9rwfvPVmcNALnP
rHW0rlHK/mTE74QtkUq7+2rThR9SmxJpFQ5cf5LEksWQZin3WMTH+dxJ2tmVLVkE
Gn3dEsjbxv1sDq2B3T8q81t5qbcfmaVuVrrOQyj1DLPQypU4JMrOVVOv2CkuQj0w
kRqAnmQ74Q1BwrgorQbk+tJpYOTpBF7phWk634EpVFY8lb4hjj0NqnWvVSmO6Ios
Bfyur0y2C4f04cmuNgqCqP3E7bYLNGPg6yDQ/g/NC4wPnBcih/DWAI221H1OKyA7
ta+u/AHhb2SKrahCWjhNslBHLRYNknjuRg56N98VMPmlzipLNx7GgfxvjN5UVYWz
wfmwWpN2Upgfa+WIVGkgec0XvA7jsz8txI1dLtIEnLeiDme29RSzF9KXWiXroGF4
vNScwB0w29eS2FuDMqYhwvYlbLgyy8CagWgTdlw4tFXy0Y7aCdTheY1cQLfKMJSC
nlRQRSxlV+qFnbDADz/Z4kaf79KWVGyi81flNbwhBpzop3vzcBt8Adjr15UmVugh
OHA3DsOwP7iBrnwBHaxzMgFnmGATGipFlO9XHawQBnyMj1VXJfVe7l3BHhTiQIaA
TK9MXc8+qx5I5Ggdx8KGLV2tQitj8EWtwSRorjN6jINoI5rMXfFjO/HiEqUlBoGf
mOY+WIm+kNF9KJvLjY8FyQuj/fdRc8YAJ+/4zaM7Ol1DGvoiuRtdkFuFUh/2rtQW
MQOuBLu70p2LvP7gryVUSkHnaSu5rZkQ8kNqCjacoR0KduXScV505c2cL5zs7CEp
MUqCtrq2z6/lwGPxlhM3ScOn7VfLXBIZHpy44ub6BwxXbfWjOv6Lbk9DE65VLf15
2L0Oi18lLHcV+pVkesmL4vDdQHZqSasbCGq3+0P1ENqlJSSXTwMo3Jvrl0ER6t/R
L06xUe8PAzun2D+ROpZ1MiDH9P3IWfdLCBLkYBCW3DzUYuRaaqVIw8aenAmsVKV3
4ij3ZruYcvhVE7wmTIMRgUA+dMZM0wczk72nyJxDr+v3snOZquX+aoaL415y/OJ5
/YBlW/MKQ73i6k1DHtiW7EQ9a8GComOVbjI1ldFLlQOh9vMAWsrZO3sC+Pgwd02y
Y9YK3ASIVbFWFCrtMSnjH3otq91GNbmF3iaZi9ON0x4vQBrKbFc9wFeQIKvr5mQG
KWwtQQT44Jcq0YeyJha3wg+R/B6tiFOWobCNRm75t0QhIvJgozWWtUHdmgt+Q1N3
YwJ/hHi5f30v20oY86dPfumqZZsRtoONUrj3AfeIzH5P4NnEvvJAn7XjLnelQiFC
TaJ7ACHf+BF6w8OOoNcZGhgEOV0mGgihu1rIzgfR5dl0FIg+Q+3wkujq/mZQvFDR
bRcMayzI3TFIJaAZ15RiN3Aq0E/qbM1G87W9ROaIs0oZ3xkZOTHmZ4pWVD4Yy0Sj
AwibagFRa0gu5KRMYcjsg6Cw2cOFMnXqW0sijAjhDhCv6wcySXxUFG6gwTmA0qO0
ve7nns9t1JmCr5jnEEBMviyjhnhoTYCDHWrcAVQ3TNG4hgmYuh7RhPF1jlBw5SEg
iVb9erVbWwS0mgS5v6o565AgV+92qOd3gR5x7rYZATX0VID1oWtR5O1vaOizUFVZ
QtaxlZ0xPQWFxlSRBXR+AtnOl+0bfOrhz1XdHfB49CIziBHvuQiH/WNsyFG+Uuez
7zLDyz3k2OL1xPniEezFF7DTr6CgZHMLo4XfRdqte7sQWswmcOHwhv3lvT0JXUAz
4wnUJV2gtwgWhpt3DWT92RSd31GpZlGWXvq6ODAXBXDTFLgN2NCtW1sEUI0YrOPb
qqAxH8F1dISv2Lm0DS7O72G+rVCDMC0O45Mf5MhsDP5mYfQSDQAuGa+cco7AjJqi
v9I4QdiRjjPApTu8CIG37JwLwRjXIqTbweFc755R4NVxMKVCQvWnkiD+PasZ2OB5
wACO9A9ILKGF9BjD5BZ3WyAomUd5c9rz4wZPf3eP+6Xemywk491ZiJL0w5VemAz7
T1RX1lx29w1ez+NWU8wYt6Wvz+LViutMrGL+t36JHgl/pSWEG5WGdl+nV0DedV/D
JWbwww5jgaNm4DrmdgvWjy0ALaryyiKUnWmAkMZAdMp0DUYS6SCtlBz6ncqV3FB+
XTD7hkrurnMzTJ9pSh1jUyngtMbxt+bObXtfaPt7AWYRSkg2HnbxBCpYWDzg2PAE
angIIkvNEjPO9ZFb4E8ZSKHbkSY4D0ICUVCTPuhLuVgi8hy6ISVZ0jz0diecnhQl
KAdtzju9wZaFE206JWzdUFpDfrBw0lkBs86cK5vvdXlu7xKqwPv2+vFdX9V6fcwl
Fj2gajwmhtFDPnMaYhUIBhbEeIh1rSKYxksUszekAHUMk/1kJYNv+3oClUQE1KEJ
rVtaEThWGsDSJLon/LA+vZmfd+pHyFO+wgKWcmCdGzywepFJ/wZlHuld6tFge8Wu
vY5eXUTNBreOW5n1vZEvOACwQN4MDnwitEJxrgK0dhbRNnUWgW8aarqKQY4trbpA
2SHswqBMUD4IrKir4OvjhCQl96ogqf4w5/rUc1jn7Y4pGvpSZN628yULneX8nm/i
u8RSG3W9DUyrCX8ibeVeFhLQb+OnZyDgyIwGu4ENXVsg6Q7CLcJ+Pvr9fjr/duaS
qvZfjlg47iFGB7i28GmBJ89o5tCvgvuXiqdB8yAzMBmSrHHLEjcfoLYoZIfKV7Ht
h/yvDZyoYeDK+IKfySzrzQeyRuqcTBrj4Oud0clWs9lHE59urXLibUZlVS5vz3jm
uTOgdPH0t8Cnf57Pfth9QxstkQBAtsy3Ws4I6vBYoSuQJUZe8NiaflkGIQFkiNxx
wpAtkr7RBznxu/hGw+wBZHWBGre62dOtUinTnhylIYabAQfzWoD/T98j/rR8NZfd
C4FrGvqBwNYq/5Hfzj2iCZD8Lt0y2f0Nktlg6LqWYbBncpqoypb9L94pSbu+Y+v/
nJo2jiZ3HFQOGVlWm6AcFkEhXMFoHWkiUF/xv8vpcZ0sZoVV/ew370aErx30NrkM
W+iFN+i7VyMd5Zhl/Kc4uY6B/Hce2xGOfZ+AIFp+KImzKn+Z8XitFTfY0ysSnoP7
9EN6asoW+e2dOpucsAfolx3QZ+Jzu2T7KWFVZfKc15FhVig0TRYpVwBUVYlVTFKw
eYFN/IAgCa4bd/kgHZf0H7GgP72j4qJI8rAuaGl1mqfrLglwsNVXEu6vu+v855FX
TthNkjz/cYRwwaQh+AodAEyYKvSJWzV0lNIiVztPQHrt+J0zeIYcgfvwnZPiCa/3
em9dThJDcGHc+CW9WvXAR6+sr61aQHUbajmFEMIiEFBtYazWZC/HGR1w5MttQiJv
smJ0x/ndANDjN1WUpwblanXH0SLB+0bEJwnl9HnY/RYYQkz3yIYz+hhLiLBU43lA
Fw0sHpfspnn1pxT9gY3OCVdZMmwFZfxeVyj8R5RzyroD9YobTVyxVqz4YwQPYHAE
xLzeXIUSZ7R2BafpoMgSaQQErbDjLLu3c+dTWjq5YZiORN6b3XCe701Pgso/PBNY
KanMWlsPlxkzwuPNi1TKxjN6GnClrFnswq3Rfrke0PDwh0WRkuNLcQsGzJvKCzp5
7uVI15WpkIeb+8pNiV/F6eb3q3tuApesBDIb+MMhjpu+DNQdvK6/F5UMTJhVmIua
zcombquh7S8WAZf9MSl14EcolOtBVTNLYyKYbEGsjcOGdtkE6pUpJkca/GEmlKyp
Ouezlzj9LCs8txCgjojmdhvHeopMYDiBktNq60yRb84jgPhF/HrSjHA0UPA3lbVO
zkbKSzvFc18Qhf7AJUbvhLqfKV5mIbHebFpe3CVSaVHMU/U6D1Q4vytWj1UxslYP
0AGaqwU+mb1hYZBR99w8SVEhvQaOsMv/FQnzy+6sp9AMBYGjKhSjQcIs6T3ynjKi
gf1xIDRpM9WqTL9O6d1vSTxUpa8BE/e1ip9MKOjred0AO7kUOlgohVeh+3rzc845
MVaXF8g4b2KuXVPXRIgunhsKg1qaPOcahe7+9I9px80Sj+jGs9g/4QUh6kSogUQk
locCWNNO8e81RVLLLBJez++6jTjPlDoHjywWjeLfAYlcGkZLAPxNAVlGzYHiYNvf
l7YpsZfV2gIp1OqBnZzOlhPM6mozseBid8eHqa7/UAO1UsHLOKUGvoCUEzgtSqRA
HXte0NCofHh5hbMDUlbxvtA7itm19tXry1n293ue/RA3uLKzsqzTpWgBX+PgcfMb
M+ujrHtrNcZQAsrNpbrGIrffrquNUK2gozAkcu/LN3Bix7KEHVvxgHeMD+NSJXGJ
YV8OPQsC0a0+0nAuTyMEbgJdygT6Kju5Agw84MQlsAA55iW7Z0Db2BxnQmPnIuo1
dZ+yUVigemv3I0R5GWa3Zy+NRb2nmecmJpDS4Pw/5Rbz7lVd1xTtu/RCSipo7ntJ
D2MMcFbtCACHLlOGS10nRJ0GiMPUMr53YOoolE1FL32+bHMmtEnycwsOjwXVSuRL
sw8jOxZWMT4bgncHhu1kSaGHNX6OuMtQeGtSOtW3HTlV03jkHm9HLBLAzI1EIl14
K6v6kAlqppts31cQ7JZqM/v6DnkpW7b/dfQYZ4+TS9NcZBlz4K/wAN11Ht717ZNi
mStZO1got90dq1+6lQnCPot/wqpDS08zTqRg/kSDut1zWygyErTAEtMqyucC6wNJ
bFJPUnpm4raUV3mqJ1yqLNX7gCjlXcrkGJcdyAkNHFGL62YGge3X7sCakALT/PDu
4cvQPZtPBZ3XBKJYnIDmf6uN43uMJ7A5LJ1MXwLaF3sAspAoMfHEPxSBfG4SZihu
KpjvGXiXf3nUQaxOBvR8SX0D+KNFbEEIzcNDUhzmdnN2Y6oy48rNCDTI2NK9WrR/
u1hbWKZOqlKz4eKWuO1GTUr9K/1xx0kAQi6sjxIIoKH46xzb11KqJ8+DlLhNv70m
zFKCy8KIrGJK7LU2whPxDPLJXM1OC5q5aJLkW4LBSpU67TVhXW3pGz+KUv9FTkTy
pRyK2mY+iQAVnerut83EGsoZrPQo1f4qGRqkAmcwyd7pX7IspUZJBiUCp0pZKPVv
RDyuCZaDGe5dXPoloyc92pWlQkiU8FjZ5lyTM+NLEJKkD/sf8/0cogPFu8A7Dcln
NUlEhvLJOfCVDkDkeMQWrXe85HOmNxEld0VCYscf3QDviOVb0umC0ey/bNUqXML2
J0dGDHTHVsr3iooT2U886pVMEg7Qp46gew5f1qkBIL6RJGfWnlXrawCtCxJmisaA
Se3R0UZs0AQw0kPiSDzbT1+tnKicYf/KgrQ4djfGMvoceaYHTvpFI4RcaaOgiKQq
H+OMTxjgcdKvq/XwGUssaw/lNv7O+HbWrbf5sJ8mgEoeW3TLYNGD1gyMCeQBT5uK
t0F+0eTIlJPjr1e1bYSbIG7Y7GeV+Fb4WT+xrSPHjJM5l97dClUDbEaCxbgC/E+1
+wqCkmAEfbTLOMHTS9z5muNzGLFUJKsQzyLx4epTccNNh+didpbHJzAN6JIXpOWd
cuPlkIWfIaK7XvE/Vxcv0tuCF535ngTf5uhMzgd1AzHwVbTGGy5WC3gH7KcIrxmw
FygPQ0IF8lmHwmf7zosedzUV+NmSOTDiT4wqj/oWHUpDZEbSMxaRvl7cs3uSQZpO
fzyLZQTG0bXztt1sSUUzXyHlTrXCs4RdshErVhp8c6o5hIIXyHHmMkis7ojE0ofA
0O+C8BQBbnXPa4l7+UETLNc1FcMBStOyH2CCpjBd4Wgfs2G7nShRbnOHBqQw22Ky
ZvRF8dfiWck3+GLzhLrrems0wjji40kUmr0tWVVC7wyHLWJSXG5qTPYiKYpoS0lz
ZVFYg5OY8L3tmKNoFPYnTuSg3gtekSUE6PB2j2pUxe5YVbKGOFjLOsSt5F4Rud14
HMlff+0jgVZXROfDabZ//+oTT9ImWA3RvLkaeGQI2cH5ht5rU3sApFxC7iv2s9gF
gsxryOfJDXr/0o4nO4WU4Ft56+ITaD9WaqdfuEOxb4NDZHemR3OloeAIYiZNDDyR
zCspVn1ht6fCs/Ti5zLOUInCKyk2J4R6B3KmRwQYJVssBM0F7ajj5ZKsE67fyfS7
IYYh5grad09cycoZiKTTb+Tcrhs0rCIzD3xspHzcM9ykEagbjwIYOCWvCG1TrGQe
TCidAThsxb7UGcdWwWYGxvOOWxaMyCmStbiNhlQvQkoEw8WSduEUI3Rxe1konoxR
EPC2Tfw5EQ590kgVDkj7p5APcYXjlaLYtHGdEZAGGz84OZEQOVaNn6gQHFqfSrcB
fqCyZtHCiJfVDpW2tOEJyIgimcmAGU0UTGv71DkNpPwzctPxGDPngrdu5nDkYXAp
Ux0QbwZsw/XeZCqIRTCYigoFUOE68ggM5ALWFdazkfawkFgNnX4oTX0jFasC65T2
l7kBKFTLp1gQYg0rfEqzTMbUP3Xi7TuMd7Wmlg6UyT1LyuPKI2SrBc6gnwCQ3KOr
c93l1Tkg1PoBMKJWMnkmHsfcQZ8HOMQzuLbXUQcmIGQDaZjKgTtNdiR1lLHpMomG
5xfk3YdZwpGB8at/WtCA9LU0YnoD15JI9hZ1KUdPBNV1VBy7VilAQI5WvLlE1f0U
VosbSVqC7Y9gn4uyiqh8+nRMeu7mPv00lWq4qgR3lrK91sh6ymxj10ahmRAMwvQy
CrvfA/D21GO6t0xHLp46gW1/063F0Giv4OPR3qKH1aaX8736+OxDoemVQtMy5a6C
GaLFa5rhvHaxLmyIuu+UcYC2u2Db8lTjFUtFpeUBQpLxgxfF1QUh0BP4JyyZddBe
QvYeQRZAoURqpe9h+JKS172uND+l90RVKX2nq8Ay74XDYBaW9WlwnyoORovssC6T
Xdhe4OvWzD9wE4jXrzuhJrEJuGYgNpxc/9A2Fme9yGdQ01HCVLGjP2pStdF4Z+RY
Ihl0QdPBaz+gK156m364AVd6N74uX5JCdcMNI+AclARiGd3oKcDdro3c1nEWolEE
Z9vaQv3ZLTXvB2N7jSo7pvT039FEzytuyTcUh9oLTiZi5yaBY3EY3Fh6KCEq3tuX
aHvSf+Ue5sWDy6pa7XbntkzB1ojRg6r60GNu3sJM4cPGNp/tUtGkBdq5kLyqpVAo
Xmv7h9VwBysxksKw7ApiZQTFlpYxOZIFJd9ZSV/uFVbEt+DwFrLKT4F1FhF++i8c
4/03V1fchhDgqnIGPkfMxS7KoEvwoJHJafjIOk53xXkUpaPnjSxIyvTxYeCst693
CpYCsYObHSFBoCvViEAYXDbrys+tJHkpTOwnZ5isvlUVis3TYcrOD5/c2w8m5ofD
c9uM/E2D21dgHehvkOQ8V9WZLksRqmnyMFB9PgpZ2YVQ95yYg7Tr/73GiLXtUFIG
753KRyCsSjmlC6xingFzQnmgIZANByOCbAiCiEaPMlr3uJ1mhTNaPAXYA55g6OvP
0ULl2MYUKOpMaVVXdFJFyprxsTj/p/BdftIMNcG1MZ823v6LL8Ox7/CVJ5xLwfsF
DyomGzV6VpffjEKhXyucusVqzluG4aU4XyG/IkXFycxrydTLoq8ki/d7W8eIAC99
uHIUwON38ckuAzEaaIid73LkOPirPN0QjvKbPN/O150cuyDX6GC8ZUMLtnue9nCk
SbG6ZkAsLQN/pFMKSBP6Jdfsss+occPMdD89T95yHzKxWuwjP4e7DSDiAzyHHdBh
zqYV8iYvC7+G9f51XpXbySRKRmQdfNNAyhVcbv1eyfROqwrebSqEz/KwluZ0J+s+
pAJu+g2KPdtOLSZHVgAiFiT6hF7thiZndYNKod19RGN6NIe9x6VRTpqWlRevT11d
T116qQeDz07ZGCMaXpNA1Id4EzvIE2QHUNZQQ30TzW5fxyee3U6DHVZ11xL3iLxP
uMpS4o6jpo4nRf4AHKphWh7btq/uqROCUiXfjxa+GUijmQ5UiUmCW7kF6kyfk1mH
6dRpEp+cs7WEUPe5dYCsnI63zaHF9JT9Hxh501gP9qqq7i2xS7F9ZR6A3Q+t2KBy
ibXj4G4vyCIEvxI9IYBszWE6pp4ad+tD16FHYmtDdjEZ0EDioDWB1hw7Cu573244
lDvYP0H+5DgmfhWu7MHhqHcxmsX/MQzL7Wz36tTKt2c8RagEvHvduH4izyKpaE6s
o9YH3ZxfNkm8K75g5pISWCt2lDsOfOw/dSiqSZ+VWwipBBcDaAX2T6pD9g8YJou0
52GsGrjdb6cvUC1xWxmEa8qRpjIL84ztF6xWOwigcNP3Li7mHSJiTXXCxVPlUPHq
Gj1tlCNsga7ULEXYH+qGAC5MwfIRA2H4WoMpCmrOydSOpxsaQxbiaeFqgdmayBUX
Qd/VTWDgoJAS9DBJMKBAUgRg4mZii2kXzcnS5lyrjvxbpJrKfM7ZGYYaOiKNme7h
5lnjPkKYVNUl6AuwE72fcN8l4GHympYTOKNBuc5X4R/AZtCwrC83noYBCDi8ppP2
A90H9Oa8E/X3LULpW+Q/sn6C1vaET43p/FRNYchr9Svjh0GvkD61qpCU+wbKrtm5
2cnco0OGZ6uetgsxJuQSJaeMswlWRwUDMSQajNq/88meqvl6HSEUzn0Joc64kPqS
bP4h8aq5mJ78+xg2IjghwwNCMfbUdTB0xPpX0IWVG3r/siSladoVm87KAbqesKTh
MfYsj64xd6LAxLf2ipBDIzRVeiXHcn99i3a1nX6lla9E/kdVVNzAHyGltr7HVjI3
lfyr93M7jtIHKrx3bYZumqfkjsyc3y6TACLRo42NCxQqTk3QuMKV9LmU3104T5x7
gt1GQC1a6QtzybFUG9d3kQpwSYY6YF8s6+HEHocZt1lGOdudpSgnfFo61+6qne6c
fh5VynFPvWQUh6eGeE+zkeXyzmDKz/ySTi3CRZ9rT5hVjuh1C5di1glKgxzVXl+8
d7y0MjJtsajYVHqTN2JsPwdG5DKe19AC1Hdr2SNL1vQnNOM+dbfFTtKVJhLv547W
EtHZrKravbCAW/OHEytK0jvBbvHmu7oDwdgEnfs0iff/cCIp9+14jwf4bg24K0Ai
Nxv9kv9hW5KYp1zQY88oSqs2OO5axRWM45Ar7D8HADM7HVihprehUQ66KWDrKK7S
HvjEWCILtqbudo7GjbbgIXZRarGwtJ9D4zardWDSzt8XZIeo0pHNzPkp2iH7kbQL
EkPAN8Xh3foxbVpckKsPAvDpWzVvgN5e3lVrW8byxmPeHXJ/GIOFJls2BYs18bcu
d6yZDgjeLDdZZs1t+cfC3tvoLmTBb82MGuSBz1uExjc1+sPEwA8nMZjknJxYXm7K
J3EfItcoKFe5hN13O5q97CqHVKx8GDiNxgfUTmVMxm9npOKyDI2Wc417aWYErfF2
9x99f+lX8s6tyhqEinGkN/mnvo/fgL7ofE4F/QSXGhED3sOJ1g5ldGGALYt021eX
7gURtjicONbnw9RZ0QCqMU2g2qVSO3XnIER6GLqWn1hc8xOBsXHmZ8Ktwyw0T3iS
nNIvGzzhImRbYpu3hrpPkpPyULYBpBjlYb9zfbKLlMk+NPBGAapmftuWO03BF4Ne
CpwKrDkONvUxYULsriiTRk+KRX/iSg6djkjbXqvVLlvr9I+bPU3PjGV3xO0yvp/h
IHSBE8tHAHS+h3CUr7krfvi2qiEL1c/JcVvbTPjPXaXxh3wKkv/A86LBSOqsbRql
Pv3irkBos834rvQ8kWW4LSox14ZriVnz4WlXuV8z/V0umahgMEaW9dUM3tREW8p5
sCbiwP9BIobVr4S02u05MdQTR00+hOv2D9wIwL860WQjJdQIWHZPbLSh4I0OlS7q
0TJG7X9lV94MZUz7hNq6efFy+LfcozWwfvuybwlIaIuFcMx6MVwCRHroSGkxoUG1
0cOJFA316N4GDItwl00UiE1j9I1F1qvRltcqIITELbWw+rii6PtVLcUG3GU5+UjQ
npYARwS4YX3H8W1AQ+Soay9qykvu4MuE07O95RZcgfE2GBfguWesx58yujSMxCfE
VVVIVRtqdnnZROON6AHT4W2444yPpBWSC2fwhubT/wxHuo5Imw8e1xsvdKD5BBjP
erJEm/N5Z16zXAtrd6ROPOchn+ZrRyRVQtRthJDUsC+UEjpDLfv3fDyS8V96wdXW
qEkjAHdESlpQqoduz3mkTtUH83mUlBF8IhFBKv9gOJdWHIj8HpmQCJlecXaW85xQ
B4UmxfRi9IzOOkeKNIIktUtz2SIHX8yjGa+3UenRnpatCuv3P6USVUPQvzCwaA4i
4HECJLBMPFzKNAo5BMhNtzy3MYaraZUGrGxq+qJmwLBylUdHa1ekJ7M0nlwp3/Hw
jB9+yZVbHY+kHfz5c9GUlzhoGgSMnwp0tjVNkpdvizssYZGIAb69op+V+s7QDrWE
uUmRWq/LFZedj1RmdI3gk/ofwf45OdVf/WzklHmRk01gz2GT3a74aQLiqOqOE/cX
g2XTHMiB6MSZG15TFOq11IwLCSy0wbLV13YHWR2D20xZYtIJACh6SP5Cguwxwv1e
eNLWWyrfi436yikYJbD8cuzRfT2+nMdUGW8lXcWrul9rJ1WkYbNYKwXTrvDnXmg/
DIRoTdftb/zsj+F6C17yIyv1yXSRxjutudtbQQtvscIAgGGpxF4pn5D1UIQGQOOU
0cAE0nbUBAlMsLMS/Zs9BeXWAFntywsaVYM519HmBXhc0+Pt8zFM6sCn3/DUdcA3
ehVkm6CMNzWdGuf/M0sCqBVeFLn7wERc4uB00IrOs95uArLBRMsJ15wAGiY30rYk
BNnY4s9CL+4hVtQDiCmrRiztN9dtZJsbu0Pvl7PmAsXfVl+2t+CiuWCnlbIb1zTz
jCUexMyoYXqPi1vXeL9FFOKNZLR3nsf22MWhxbFdEEYpPx86uAg6FYJF3EoznY9U
1WFwL4QHGGvYiLLyj3YsifCKqtKsk4jV5y0/vCuVjx4Mmt+vmigip7x6P7DDNns0
jIy3d4abnmfwGT1INBamh4b9Bwd7S0yDd8KolD0lf5Jr11P3qB36g/gm+ZUUlbuJ
ZhZFHhaa9mvDnmbODPYug2iaVUv+e6KfsL0NxiD+e5IaLCCWntboXtpnIxxD5xTV
wDmxsna3Cs/QLGuY+I2TmlhP0njxhyGIww9yRhyS2Lve8TlXMaQeFWF8CDaSL2LQ
ocEnFUHRU2Fl5TmTmyX5LgAkqfaM51TbmEtB/TOFOOqVk0v4w9s+IZtkr7C5b3Cs
PqwqFC6007NxtA8hYL/UFCt1l/9hG1Z6IY0st+IMxb/fQwW+4kXhUmpm3XUfvzBQ
wI/r9bX9SQEHwlKgrCZAtuZ0N5/2pIEb9G0usvyBI5btyYKwHEi2PQVRcRrefdCr
wvBquWJuLBH9mlg1ZLzryc/MiaXhFzBwLH+gMNhhVk/lZSRVCw7qs8UyJ+xaH2sI
gY7Pgolf+8CISbAFInXYJzvBxr6uL5isxjHrlb0fnwlJS/yB4/cssSgHqIwGRL/m
Vf9SdDEd6qWhxXQj7Sg7FRVR48TgSfmM6gpx1t96ar1jDiV+/64pqLkVtYXOoCpa
X5PtHiwYPwkfJaPdMPgW5NEW+eDY+mXodnpdoG6v7qnnd7d5jBSQ5VeYUAb2oXNM
1HYZoC7zuwmNLecjgxl/6Os4HBtrBRVOhDOh2w+HtId+lP6B1RL/dj+8xhPoBlvJ
YijKcINivnaQ56FFyBXO3vlieIcVoP04aJtCfP3rpZMq9Sis3BkEfYpzYp/JYqWN
klTpsN0dnStf6TPwySoB2C0s/e7Moj+y52h9y4aVuHzQKFFOEGS4kGH2SXW8dxIg
tknuNsXYicqLTqQ+xWd9KzeaVCqqKvO/ZqVQH4BJhE+MLBnT8eiFwvLbG4zbdeqe
3YYFgtsPe56NV6VMY6+DnE/DTk+rynmVGxygndw37gkxLcRaBM81qZCnOsNpRbhx
gqiIOmDRdQIM1EvXy4HZ5m6IilbV5gvwp5QRZGRsE00XOTq4q3C+J3lUUf/192L3
X1O8OruUgSlPKuOXxYXjcpboUt5XjgcA2kpLZ6/YNMr9HEriGLyVJ1CnctYAjCDc
gm9WJR8S0uw5XKSAW83LXj9hpI27XD2zJ6oy9g7uCac2C9c0SVMjASwWZapEOeR9
Ufc6YiQFylUMGSybzqSKYPR5vgLS50JGq0QVFGy7EWADmXJApCRdTmcy7sC7mKVR
wkqwLK6LRaHu+oc9V/4N3MK1xc6AXZJkeJbJdXNcqlntyUOYrK3eNSKp0sqUiZq9
1HmnE92hTCBZOX/YCaGFFHtN4viJ3zIo7XVVkmfimLkuCDsxYZ+VN2NwgPHZvscQ
Qw9sbhmH003eOJwb/ukeX2EQgy1zHXvMIDiru2VVziGWv2ZF21N3zDBD9kaziFoA
iFYN7rpVpb52UukAC07qRh2Go04i+7fB/Duf1gArIQnpHWZ4lHKX3W9rUyCl89su
c/KbmvRRPsLqHN+JGuzl4oPrM6rKXXNyKkK4mlS3ch4BSFQZZiXPwotUHMxUWLMk
GwYkkzYl6WYAAWfscB6Y7/tC2UvcHmPQyXNBySm/V48FT0Yp9p7kqCmdQmpsRZBo
9qQLfflhiiE1WTAelWZQn0zeybjOgTgdJ+I6jTgtPFLhRFjG22V2w2TpB8C8cLY3
NW/0kTB7xsmyvaZaI5/2OKvWtTViHCbSolUuNdmmCrY4EykYO6cdcvSu5xXTZLkx
xwxsTPugrqE7qYTnsVfUj5w8UmEs3whEgtpO9k8ta9UCo5FGRq/CrahrtyxGbr70
PKfzwEYqoxzm9878rd+AwKYMm2UYyIaDh5hnwfuAzHcihb+iOzdGZQH4fzG0b28h
ndVHMYRlW4QCAx5fDrPyWF8q9iWd+O1qycs3tQ/g0+1mTBZfS/1XQoS8Csd+lbon
q4SLr1NkyAtdMu2DT7hJXBSMGXHrkYGIttVH/v5SNszw25WIgZhh/GFnOE0B+HDe
cHLzPjohqEQegyxvlfnm5TWh0Ay5mpumyrhDOQsSFaOSfififmPDRk+oN0guK51W
Kf2wg+AFdTmb5WLIZOiQrK9zI6U25Ofh02yrxXVykglyFMljA75UAvi6jiVJHW8q
dZD7dFRcRWml/KDIuKveiYddA9Fz9c8OLKkaSvGqocBZpHUrPevI+k9lv8DD79fa
wWw4fMvcuXSBj9Vqyw7cGUAd6EzGQlmWOYlNNA2jIUfuePczu7duNMh0PtsJJscT
y3qZq+/IwDkPehSGNMrS6aZ5/eICTkPHSUxs/27FK5CP7yeZI97EU13G9A9P2UIb
OrypO2oFKJ6vaVt5S3yPmzLe8QnXZJmM8tPZzJAM9guJSNDGLXP6RGbW9b1QcMID
/ykLH1Y5NZWKiFesnMAm3dzl1H/CRQ+NZ4KvFH3INvQsw/yUeOIJuoYLL2eADPwu
CzSYqzBLRQKBc6ruvwO3iubh6ay7VOJCPE7zHQo5WOC+QYfK+ei6EaTUe0ECgONC
LJhOlsRb3XAqb4hcvCHKS4MDiQ0OmrUTpK4liSkBXc8fIWkhHFtQJDI+JYh4nQrL
3kAolulylDkmlXWwZM5BRFFAqWFxb7ZREvby35NN7Zg6sGW5AqEc3o9irYbVZMCF
32G+DFqSPKMfUjJt2kYEFFvYO5AYNbMMbBRpprpfmTmBoYqUleHBeepMhwbY6ABp
mf0/sPalt+QX9L69eUqFk4xb1fALhQFa25wa95e/yp0ThtXASAUG/qbpWqrFhSDU
VxlYBSajEJZAHI9BhXVtzi1IbV/tvHFMidiMiUH9ehfodwmBE0exg2UufakAh5X1
mPKmLNAwAb89aN5C3CirmiB4Ohs9I0l+YaPYVKoV3u5Pr0xB6XnBZyIkrPWVbl6e
1eK2N9sDUANqbeKe/yi+gNEaGXf5KjuNkFOm32OzcUYO35qMM85bTgG9UFkpcklH
sCsK0G/kSelHkp4xzmXllm5joR/ymwpNQ6W9zrFKwQfAVJGvIvWXK0RueTLvRMq1
et9KD5eLizG2ut8agki5bwKWWrVVYjTddbJcsW+FiElIsZEj3cTj5ouQZ/eY2eqI
VXsU4RdbYOJgdJe9ysRp4Zesl0LCj1r7FMGYA/rYKULybQcwi5imdynJB1c5QKc3
3uOz1zisB/gx7HYKGOIDCy7v6I3efZJLMZ3Of7uq8/sPa9fx7lgWDV0wQ6/aBpO/
DcJBOvKf5d4Tiz9Cc/jsU9HOcwRip645ZovQBBm2rV+rMWnw3ChRi3RiExLY7aFJ
J0KdFePJjk2rTMZJah1nc4xZivvyfKX+Vrf3THG1COaHx6+iWw2TvscOHG5nPr4N
DGm+h1Dq0J9m9q5U5LJgcyzLYrjwjdbjDeOZ5GiZGvA/s75Mccc5pb6MGZ9GJpdE
nO5fBd43eBJJXN2HogRuVonWkVsyYR//bds/uEfnvzQp1cA5e2qKHnqKEZ2tzx2N
HYlug7JgiljWo/JBgAd6Q8FqVS92l1BuE5e+iLWSwFVtcQsSRszPDzGCsOv6l6ou
s1lTbhytJlILJLZw2FexlBl7I4aGCbG45wb66opiLAT/UvkWyDL5IHkM9l8w29ss
vfpFpWqkCyrq/m+/ZV1ML4s/xr72snw10qZMmfmFt8gyMXgtNigoFBSfXC9NSsPS
MbszsTDbVTw6jKb7uTwz/LhrJadhFQYS25o7sw/P1ASwBSGZme43aCbk5kEN4g+E
Q50BkuaQOp5Ntov9XrESXbVRW9t3RJPPGYNFx4P307K/g9GXxCMWUl8Xag2p+j5Q
2LDeQ0nJ/FnJvK3vgxLaaA5abVr3i25EM4XwLc59G/gVodNK7ANAb3VTncmyT1eJ
toTfC0aswnzHYC2fge2fssVriVxual025evaCUWV9rvs1JM69YUvZEM28HkagkaA
FPBPAMgue4BG6hRTUKQV4w1WSedOPDGRe3ywVUoIsAfezBmUPA013Y4YtCDxqZKR
B6vURUhR1I01PS9fAUsfz8u4b1d8WDyCiQoaNTctvNWQ7dEOGv7TeDyoqBV/te2m
DFAElie3VP7CmccVEYUXC2LptB4VkiLtLkAn5eZ39BwvY9GMj/M6xYh81WDSNMqK
cIZjiUXJxLYzp4xT9mc0mprYjWZTqGlhfHdrz7We80vRJAVGRDuUvqkWVVKoJB3Y
10Bdik5UzjnoVZ08wKkd7vqpPzDdc9W+xKObL/q/xIj0d/70yxL/Ted1KBqt8arc
FbgwxIzEyhw68f+4D1vnB7Y75cSFApPGx5sDCxPDBt854tsm3uocqFodxa7qUAan
wYdpYRrtDIvwQ9JFPt9CO83rbiFyw2aqqiU0IsM1lJSzIHCC85pJK3hPUnVbr2lw
g4VDlUi39OaPqK+FdHXAqzpgEyaz2TTeTigp6bIcpvLGvpz8hAnvk3qu2Dwsr16D
7d/xLlaFhdqiXh9mfDsQeXnSPiFBDVr0payNBOQJeUXDMB/SzuxZApNRFe2lqYT6
ealby4qCUCx8wiaYx8X8k04lwrEbsraNdNjp2GofUtTnaY8BpJKPAT1eoqxCK0cQ
VhzspO6svoImmWBUUidTOdmA27QleGffPImJDziBzS4PiVWyNCLDqagDUe4Kpm91
KzQ6H9niAgTGOKt7azdsoedBmoKk4julgaIJX8kHSs8HF5dVNOVbJj0tKwY79O+f
gBKgGcYOYTVR/JNczH8jRUAWI6VtfqlxLTKMKPHAgd+Q7/8NhCCt43oR9IppQMYf
/838576SumTHzt2y9YE7xs07Wdzo62/JgtcTq/v0/JGPpvGp26QTRbZR0+x0Z5Cj
a9aejXIBm7+Yftq4s+RQrDi6g4x0EwuSvgZzEu+V/2UgtW1q2TlJhPFlJx6AhjlW
aH0TzY+UnJJ7TkKfZQWAnZdoxgLmlI5jWrDzI6CVg7HAjgcmUCsXqrBJcHO4iC1E
X94CAGvzlhwdVEkCYch/BP6+6A0sG5vzGioQ8PFKfFoiFX4sFPBcTBq/9Bt7B6E2
XnPBAhnHq0ZgJV6fUo5vBsngOjbs1lxp+cD6wJS+EIkx4MORa7JUgK3XWiRvD63D
kZK3zlus7yWcTo3hs1O5/j6YBU084VjABXawtoCplKKLaTdMGXFNWs9p7dCzS8l3
DInRe2ZaB0ZkAb46yWLnUmSqDFwf4v+NGBUh4Hxx/pEQdtOCt8XXRzS5lWJvL4Vj
THYfoJDbmB7rpZP95e3dqqrAEQ2muyiA3dN/wLtM6yGpn9/hTwtmiiAqitxKfjUT
XmwexoIMUL+WsCql1azCgcQCVqdVKhSrrc10xLSU4apXLDOWsQNeT1vbqhxCenAl
/r2Hsxwnx/Ug2anVBIQtQe96oWULCbqDje+DWqU1F/c07XNl/aRPdPNyUGNEs/95
VE7HgXNm7is5ZGLiY8PGgAta9888EZi2sEbujQ7wHqftXHnpiCWRxIraaRuE3DH+
cOXoUrFhHEmEi1OyqOG/wEn/ADzJ3RT19tEjO51DKFd00R6d+ctTmvJanMn3HM1k
9FxTXYiXTteSHny6wxQ5byOUoI7L3fe9svoiu6kn29LtPKfyqf8lVbzrNXKLsSCs
YcXMIknBTsisJ3/HuDmn9PhEr8IuGMszGBEWvQ4YttoTCv7LgX2gygO3iQnMR5z8
naW526TIQq5r8uU1bOqsdf2JkWcMkXV9fyk8VlrBNU6foJ1tGuDjinWGT1yvB0+v
qL6mArWiWy0qC8f1AG1EGftJNoWc6YWelPQwBbLmKEMtSkJu2fyt0T41iUfXwjjA
PCmlzT0XCSrhCA2qcsbZyzuLFU3UQzDttwiHNOijIMruEvUo8pVTJo/TGni/2R4U
HQ6QGft7fcKeK2eWNQYmdDIcUUm8uyQkD3bib+o+DvneArtVm30BNrmCGCUhf761
HaXQ/ff4+33TzHSNJmy+svrU7/3aXWoNQ/DlP7NNobqSPRqYtm62CwDdwUpFKOtN
63yrwgkBnwxxw2OtPEDbkxEIhbM8w7zQ+5q3IhHJCiE+d4I5Gzqozc5KlHxv/2Xc
FSe3Q4rZaAf6sh0A6XIuGiuqte3Bxh8A3bT5Ykgvp4qshlZjH0VGc581zyZIeR1A
ngbXyNtJzO0XmZmT2IEVqsyQpVZu8SNQAjAYM5kPhpYNTcazyBJGFQh6z6pw7T6J
XgmjmACapAH6oQ9EcTxaUgwecc/aKdOzR37OC4ywtHl/Y8zFAqCFToHzi07Irahv
mU0BEXH9TidNhbTmFKwmgAiNFubUDRKXBfPnC0cF5xzNoQpDSsYPKGJR/4gSfcwT
1Gq2OsF11R6Px0eRGgOa4wonKQoMEgKofSo632DJWw31fMdRbeNMirYQTk42KgCQ
q6aZdO7em4blQh/kWN+TmoYg45UCerc2ZjwfGs6ncCXl+er+dNeqwSxoWmTWOzxP
NjWIb0h6EG6IW+cPRPTHuRqCAk75/pESOfnmPbBo+sUzglhVxLtNEeAIFp1Qkb8T
Bf873uoCamQ9t2KuiKuK1THRv0sm9us1bnKptIimfGqr6+YErY3NkOH2nEELVxJ+
eL4FTLT1mQwEd+nm4B8BYxTKu21DtbqIuVH3zc1+LU/P2nQWD8iuEwqFUnyMGERB
+Vz/RstNOXCrDfafrckdwyz8kjD36TPRVMs/4YW8SSNGoeC428d0V04++PJLvAd0
Zbmv0bPI6M97aiOd/JwFQaDI4FcqUJoUmgByR38OaXYMOEOPPUC866+vE8tRMjrO
Mxn8FfqIw9AHCcxQy9zMtpq+KPUFImEMTOU1q11ybupXBTWBcF4nPoxBCNXqqRUf
LGe1PQlcj/Yii/IqwTlmJ0jgdOEmaIK85yfw5qJbG9Ro/pyYFPMJxpNh8VWC6FCx
mveuMkVE/4DtFoQFjRuImgCFyrdal+mrLWHwfpFky2gPWNGdDCETzDO6qElMd4Iw
OoTmAH51DOax5GbZCfCuHfC7Id5RaI2d+Va6v3lwyt+6WpJWMi5YbMcnXVkwzS3i
T9IV6Ld6GnGuq8GxirDyb+hZbWlmseWV1bBgEFIqZA6o+TSlf4cngmxyJjV5IPc6
Rv2tyXTnCOOIocBppwsTAsCF2PXP2rDH+5xds0xiPG1ymoccq++/qeNkQ4CbcBwO
IFkFymw98rEdLGVgGO7YDskHRd8qbE/j6cO1rNlduPwmO5mSNRYTtn39hmUmLLq7
9V1c6m2c2vuifxRzX45UbBKV1WZrDwgWYW8JYmJygx9EdBw+AZl1kXQsqQ95wFW1
ehYniD4MEl3fz7HeuET7M0z7c26NFnhSWnKlKniqx0dEPqQW9Wp1DUlPceG8D2Xz
rtJP7huAhPHV7GeIYy7CVYCed9tweMAqCGBVXELlQZ/fCzIDeCdiuSllrUJMzHqP
GoGyJQ1yqZBgm9rpomapbKUUYA2qHUtl1kzyZjeMfu4I7toyesZoAdSkJ1pKAfRE
O7xdFEfw/NFEKZMMo4PvlUZHBTjAUyaOuL7oOxxoc+SetjT1GApP8D7gw77a3Meh
pYek+AejamO6tBK4ug3maXmDIO99JJIyY7M5soFR383RkfffgW7t5mqtKn8IOCao
lxVIZwL3iufLaqVPnR8m04spnI7uk42DXPwPD8K6HQWlw0mbv1Mj7PwefzkCxtwR
1+AzoBj3V/GOypgtE3qvnaYyRiDA8CflO3Te7ytK1CgZhSecMKcJ6dsvcWm78+l9
FNPUJhtCZD0a5y3pXHO3MxEeIlfctN5wCYTz1WMBtLMsOJfPcCF/xLha2OEA3b5h
KwFb3e1oQQP4PJcK3z1V6FQUhl0r2ggfL5SeOZ5Yx1JNDgbYbM/CGVZjp1SN8iVY
A4cZwBDle1PpHERHwogk3pnn0/zmR4iFVMo/y6tMGH3HX/Ht/WHyjb3AR5Fvrq+d
gUDT9U7T3T1oDLxOUC4xyCeLM1BY5z5C7Wg9pZxg7z6VMso1JoKYP/Y3YacayJ9U
w1bBntA3QWFSS6FwPkR1LcorUHrHIQpYTMk0XRVoD00/rUF6Di5B+yb0CYLKa1+v
Wq2ZXtq0Gmc3hcLZq93YYE9o2bAhBqARsZWylOjdQyfLeVRbkPPdczyg0774IuNh
0qV0FS3jknDnVhKFLLVXaUpCd7Rf3PFNrvr+xoSlZGs3zEyuX5nGZZmXPCUCfm4K
Thn2aNIRXO9Biwlxh+EiLwwWWdKqM04waNK6wbwgPsb3z6NDn91jyV/XG3sKYKCc
r0CJC1PzFsGnm0CIUMLe0ee+O/S47qoEM91DY/s/15keo6FwY/n3CMeuWdCRULWf
W8C5YwBb4wXYkpTnS9LQSaerYazNy5N9Pf395nalggHdADlRRP9MiwYm0OTL+AJ7
IrXM/8nJxmbSSRPoIj84q7Zvo6D/a1AAmzc3xdrzvi9hDsDwBT+MsOpX2pFmFWzL
s7FNVqyoyTbHVVpTXAaYsnl3xx7INnSfuXWSKrX5GKiECBlD4VXWfEBZN9OIbXZb
y0OelS27Dp5/WGy3dqrgPXFcWLiCOk9ZYTofN21aOEgYsKbOlHrfPcOFCofaqhlL
AqLoaTygeZIIKkZ/aRR0G4hgssdHJ4Oki8WGrnA0yCg137eESXvp5ez+Kr2zcERm
o+Od7oasSw79Ivv7u0PbCce3mWwCtNK1XsGZ21QyY/BVuOPz4oGfPPmG3/riwWzj
JJEaO7nPyKLrmOgm+6eL2z6o79oiMokc1vkb5W09AXkRugnurVk9Ns8fmegACv0Y
Pd7tAqpveUIr/py/TnE2g8nPPcJXT+QV6dVkT61AtBh1M7wa3doqzjF78T4hfigk
hN22/a1RLSr2yqjI178YTKCh7c0CUuqw6bKcvB9fjxZi1GQiC0MekTbuGfDtbjVx
fwc87hJyTHC/R9+1P0L6AbnXvBcfpTPlpi+etiOuT17TaI29soYo8W4+lEIrnkAD
fiGjcGja2EX3eHKB7c5ZjOKaxSqZYPswEegNHIkUHhVtVZThy/SLTfuSA+BtIZ3y
4ZNjRFIcZ9yplZ8JTie51WJQqDcisGIfI1uUUzlLnGeOh+0KUrGi6v5gte+pEC1r
/enGE8UhVJb4DkJNVnvxnbcuvQp/ktu7fBGbK/U+MeGwiurF9D7GUTZhxzizNO7v
sOp91R1ttZ2WVUvo5aIpNTJqNybH6JP/0vWg9sww7LNCnUglM/iQc1hecu2+S23k
fZrgO2+JBZSgIR8B/9D3lsC7s6Z8nu6N8pCcqA3hpyD5LBb80diNp2FPayuLDoTn
9mgfs59DA9/lEFD0KiSkTU3v3DnkcWrSlZZjZSykJxc83G3ZBgz92GiseXYDZ8bV
6c6vEzOVDACTvYBVSDCMCowzUn3yeiK0vL0ZTHK8chNycn3e8WgbQtCH6S9WZacm
vvC8KDAyyRpJRs4bN5e6LAty/1l8gZy7ukiuAJa/TEXHF+Oc4GOAUIJz0LZe0zVR
uym9scsbwr4KcnbHfjaQbJ7Y+TrpxPRybEEHTcU+nvD/Ac3J6kmlJSW3eGIn4A8f
QOMtu1aSTf9dUVFqg6aIKzgzrIXMklwEAqRww2xdN4mgV/VMalkKKMCCbwowNawO
/F10FFD4dwTk80s7/1vHkIZzNkKr7zUP5+8FtaVdNl9B7E82d2Mg5L4/yRu90/SF
LdUQdzEbK7F1wJEWr1uBEhJy6/2CC16shl7CamBaXwDDrLgriy3aUPiLWAqDCQUJ
4sxu6E4n+J2cVR5RWNMXA72KxfB6Q/PAlc02SzebqsaoiJVgdlH9Cld87aW2rOK8
9XY1V4H79BaM5WTPi5rwRa2gS6K3VTSoPcXntOijDD/Rm5H9jGJxE8TxtlY4bA2B
CA5M1TdfgZuoxO+s9cgUssS9QyQbznvnLLsEIo+F4foUNh1/Agk1nGV//C42ig2s
sZ/70yrwn+f25oR4V0syMWz0LaxB87sNcoG7VHZQr66Qv37YKXYbTJ6UoT6RAt/l
oc8GYh6V7gjroOLB7CIlUlAqi2+jXXk93PVihHmojC4gnRxW3unBG9LnDtUqdukq
w+2J/f5/uY3GzK/JwfY3x+hzFl3jzIAiT9yWz7pqO3928E8B7w4qg/e6k6c4DbQ7
EZcH5H2omR5wEjfVU5f3QS7XRZHc2F6iU1+OkK8pjGVF+RwkQWn8EGiJi8gOIphV
YefmNJlEHT1pchQNnq/G+xJMzByVuBJOntJZkcfpa3QNKVeuUHCNTG2cRXmFGOvn
i9VYG0VK9duigiwfM7iu7RHod2QeS50T4o/JG1B0w/SSEg+m3Bzey8JKfH6+Tqtt
6zMVdv1iLvcwCSNZ7ItWMgI63Go8O3dpWGMa/8rdFsw6jFqro+p3xRd6dvB+KuDt
CdllBfuBdWpSwXTYRwHiweqsCt3QiebVvIfx+Q556o+1jNRrMEiA/UsGYx2MrOc2
XY/2BgjTETE6kE+hiJk9t1pGz5eRZW9+lPBlKUzRMpyHsGgI3CzBMGkn/O9RWPSe
zBjsBpCcJuNzji6xYe+D0aUHafw88E9iXeRWyfnxWU9vFF47fjHtoIY/C3eK2mtK
yuKdojqe7NgK3XIAWVriW3GX7IwzsXN3w3bbFbYVgxR51Iy29qXRGLHda8ixbGxP
YsQ3ZGAaHecGL7zDTK2zQeCsVOCCezkaQz1+VNaUt57Reah+xyhmN3+TD8grbcc5
/XFSdg/StkVwszPoG3wgF91+r8UMgqrMW8gVLi+Asyhp4JRNLiUz6xXq+FPwSvev
xDBOpoF+RWvpQjHu/irAbzDLVYqg01uRreg1h9f2g0/iyuu952u7Rzq4+hwqvsp/
k3rZWtHZOcyLKyR3ix2AHNKxIZjmVWO+FFVntj2kXwBV78lA4scAfb0/1YPIl8Db
sl5Z6m8ZyLLowl0RErR1tS/YiU6kH9ZiSRWOOX9jpokAvAzyv9f50U8d/uvVmXIn
47JR6mHsa9CPiAmTvhCIKgEOi2qaTV6CJ5VzWav5yB1d+8edWu5f4zzjlncI+/fU
TiFlJsxBfW+FQixfv5o7kJ402Gc1N/O6Sn8/s+m0xVKCDvU/Tbqbos7S5BtdiNHx
jze6BZqbGkbXK8SSmdr8CihZU1EF1dl7WrSX9qKtk/67osYlisq1zSPSO0Hiovyn
+5ptx5i72b9727seobfQLd4JvZQPz93m/i325Iv44a88PIkIMBPpod2zIo69oh1q
l7XtsEPUq5NTYbJW9tZjbLveJYAB9oXVkLfIoStcKCKH8ysRxjGVxoMmBe879gFG
JLQ3OJ5e7yBH10Z5sD5Yy5GbQ9tq6c8KWaEDkf1RNx886idmQLPEpz0WFPuGEGkS
ElgxRP2DN3iZ/FRGcvt0u0MIT7e22NybKh5T+otd+SZ7Wy+A2zPVJ0a0z7HxtNi+
ockmUzGlaQVUEZYlp912An66oZe0i4eJkzi2mNgZwGSC4bBGwfmTZWaeVMLmEuJ3
rBDVsclKSyqYXFfWL/ITHQZ9ul3y6TwukPqL//gyJDqar5PYE7fXkR3n204qkLxT
zeKb+ve2QmIOKym0epQ6bNG5Jco6S6vZAp6yMxcRfgOrq5yfHtGQkCRMzP9Mg0VQ
XgY4vqp42gQ4rkf6YKqLk3kjKB8UZrqh5kqeCC30z6Cj7ZazQxJhFfMu9yzIS6QJ
31KC35LHNZOrsvBlddisHPvFrtgx3YWEbdsEOdfwg4MDPz8hd8dGj8RRTbDbacWE
m/T9ijA69I+koslviAews1NeQ6QIxhCVR0Yb2VBVhsDxOBwb/Lv4CtEh0LDxCWSb
5NM7uWxZpvIMwOVI16BeJ7Rq9QCPzXkzJJyvaBUdIaD8aFcpjWkzbPki83gFcu8A
R0cLXwWnWQZ5XHLJCOYhURNdRaRtgGyNjJTg6H/ixqb4xSviPH671g/0gz6DCzsv
Zy430EBZkIc8wAxiq7vGUF1CESBg5BFOmS3alh6VZnU=
`pragma protect end_protected
