// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jpI4a8HSEflfKyfHG4clA5EnSNHS4RhQv9kGaAY4ebtRs4/ULs5Q3e+AUZXdFaGrWYeorTWRouBe
UTAnTuOwVe360Qu6fjWOsT/iRUY3HfdWPYy+QbQdljrjgWfhvQ3CfulmpyctTu73BOz2vlw13yYS
5UNqex0kMRWZxjqFcKC5H4BbZk7joSOV7ToxKjddgchEAKrT4sn+4C06LxzQydH6iKazhpZJVKlm
HrBdAHOo6iXn2ydvsbRDE3wLvOcv+eli7l7MinRTyG9OFICoulv1y1MNZjOxU3rvNpRAbnnmP091
1kKzoDkYVoT+4/qhmeLbHAMvm3yRA4WAnPt6UQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
0jRqTH/T/VsPmyisPZ1+WjnluhTQSlkq26UrFPhfTTwlTHPd+aq78iOUC2Ty3aIhBJrRDlGNdYAA
dXEayZdQLfaB01ab0N5SKKUHVFUsWHStlIafyTGjgl92kf2OytokoaKcaUVkgFSiacYCkdG1+slc
TuXfnRPdA9yFAWzdKghhJif92E/Pu+Pwa+WkxlEDCNwL40HKCWCkcynPpvKxM0RTrK1gWhvFA3Ip
OmulmSGrZthVx+7fptn4r3wtGKsJptEJUqhZ5N5R37IhGnDmhXD8f+Eqs26jEI9SJbMhgseNQpZ/
QcExWE1sYw7FGyusStMYTEa3jT6JzHEqv1boZnpQvCqBSGLK4KxiYVs+fCHUtQ8gncsapE3igeoZ
wjsarinyLY2aptcr3kf9RJ6eHAZd/PLK8K6ntS4gbCNONKiOefXIFFeZPjxHR+7Z4U36LLGyWXpX
oejIOz1qKyoDT4sR2fgUS0YMPN9OIVf6AHPWHnGki0w7yudQDG3MbRFF067LI8tm5pbEwZRAMzVT
lxh/MGi7aOnpiAG1MdZOcb30zAFYN/jLqUWRhVRQ29szutftELqSsL9SIoxGJnWAY/Jcu8j0M8bo
Da4Yzrv3rraIqNW6KdKrSi2oLxrZrwTSlc5qJWwkU7VW6yVtpwgOHmGZJ4hpb2XNhhPQtf/GKzvT
eerBSmQ+lG4a7N6lqpLvNRF1eRPqcihYD8GDj6Pz05nSvAOY95zMb5VCYRqK96xRBqrNsE+oHJxn
V06fPpPs0QWBgiyl+RByIQ2xE8Ou6JQjuueorXd2e6pffbrnqY2EMZvohC30m1RGujNp3qIe77cH
TxF4ZMkRrI+PtKcF5Z7ABSWeGkdV6uhnnbUEkyd4MjrQYwILfXVeugG9FTDIVay07ntH4h3n4D+M
z3a0IkEY81wgET9Rmo9S173OCJyjD0dBrPjgqgFD2HMScuPmZ0Qe0at9qW3xHjvntABMKNVdmWal
4rDO1Rz/lvzWPQCysKSEjnl+Hed/ef9OEpMHUPQsg6TNfpHyZXH4ZPx1IgG3TTBSqfsto9ahhHGs
Fi2IqNfICgk8anLNvBBx0VGL18vtCCTT/2WK5ddxI79Xpil5R8EkWGhDmw7wuF4BQz25TFvbCJ/h
dVQB4XApnLFz2+xZ4iPLr3SuGQrnIkNcncCgdYRjqMDM5MYaMqMZKQHRNn32OCQDzKzb6oXqnWKS
RvpuewovJHLo8JtE9cu9AP5pAoZY+qB+/zPw35/N8tYByJtZBdcuagitUXZWi1twcDRQDUboI42H
1suDALZAdtoGBb1QduG2QGzHPypW6+CaUx0axdKH3bjYsekHioU7yWseZ/2CsUuTVP2gVYDPaioc
wvPeiCMcato8fgCMg+EHMIfOXAtn1qWMmtCx/pNQjwOmO1Y+lnwW6cCVBexml8yimxgRlwwnHkso
MnGWE7oAhz8RjCtyJxNWMKLTlgGTNuGqKmhJp07JXgCDmMCuINj1WlY/lFsmfsCjYEJgRouA5l0O
dg3WabGD5dpZ852BoX4fbmRZ8o6XU/S9iai137B1qTVT71aipGiskWvtNFukX9MlUU9ZMkupfBDo
PW3HtsMt6CjwHpTxWuhfZmilzjyLncIJS2TTAsS09kqolAMRsdfElkooJVVMVLtoyc8dR4Xw1mVR
NQJGrbcioUUxGsypgw9VNgy7DMi/ZqLtEl9hGvifTdWzz1F5ScObI6WLbAgM+V1bdTY44fkM6ycK
e+ZMCSayIBpkehGuHt+mDGph5kK2IalD/VCKzT8gABoW/FMroDXZHqpXmtuiGXntlMCT+vw8Lrgq
KxGmKBIutiPRq+upiiLWpj+02VpxUkZvC9cID5XKcjSVK9zocBPesuCYRW8DRS/7Oi/dkvu0yu4A
olD3mcczjCGe81K9qFj2vJejO1DdJ0/dFlvzQ2VNQAXu7+KqZjfx5GwPdH43cXEX605ssmbeb2Td
ZTv9W1Z+wTrb0KLluKuBxz/9apEuoe5P5GW6peWeNAlRjPw2Gv9QQEYU8u3RzsMkYatFA7AKbOVi
Ue97K9XApzTYPt+S1Xw5cgoVr2FBe5Z0QOCEwLugzHmlg/gh0RXWwfzrt+v+5ca5jCXrVVuX6IYK
+8qBAO7mPHwoSHlLP1vpWv1wDT1+tE6OjXZ025FGVYSIt/AwHcWv5iMk/xNxdChqFWb3tPZkapVe
p7Y2whiqsTk/iT+75BRbsJbF6fwCroMpkKtYiuifuiAIYODNaOFUi0qaHuAc9T3BtPMsvC+Gyb7s
Y79BOOhltRpu5JthnhjboTTfW10/iydUEsFK5D9d3BqEYDhZfOt9fS+lmYnDJYIqfjZRw5z4T8Rz
02tfS5IUTlcgKwhRqC1xgHneN9d5QxHXZQgW/z8jUd/FdjpV73qu6JQm/qxLsxTGOPDNzgdqQOjF
AkvYAHA6mTdhi4TNKNJIkuBQA4wsY5PAXhKxeMBu4FX/xwQxdhkBouzNck4E9Dp9OYDA1Yp0RS+v
bQfkBlHqE6fvM8EfrAxU2ZoPQKmV3FyK2hB5CCn+CWuW+yJizZuB8FigK/2fBUfNioI+iYuKUPYA
1AYq+wNgymE3s1xbdg/7kaFE0ab1q6Vk6H3XcIF7pzDKwTpjJngQmi449m24FOfwEWFCMmdfYWJ+
vHC15/f+C4mAx5JtwAjCqRbt+B5b0AdG4EsfF37VqQd/YYxlf5XZRIIyn1Uy3MJDt+Vyjspe1WLz
/9dqERaJALa3er9Cr9dSzSRlDsazcZMye1BZpFrwYoRC7XYQWpupmg50jL5d96ZnLHpS6Y9myt3T
g3ZXX9QFU9nC7X3Fq7QuVwge7WLp3X29FEHTNdSxmg2j2m3lXNV+FWhl/4NgCYqYj/UR5Y/frn/t
di+goykN+kEhXwoyZa8QfWqIbVI1kimrWBsPTMsV6NdclZVDVOmY6dUCnDAJ4JJqYe0MQv5w+vtm
jgJA1BTxZSYOtIjpPMv7l6G8y2AhKwgdwpuL0bAmodBylzGqBnWml+Saqg3sLTDdykc0ZoZMcLFY
fcG/+PChfewcM30l+6mYrEQ9LetGIxYblCN2du/HB+bwEOG2VXtUXBMBZYv15aGmOUY8NlKu1RRJ
xQwLG4HEs9GmvCzmmgXFlp0KJKKbU3RyhH9PM6piymiRLZZxoKQOumPC/C1hxt+qMshoRbzRUL/f
zKQ24e376MGSAvoKlBD7LLlJ+AaMm5Pn+zKR28XlnTq7qSzXhJl3PLraiSIlO5Rnn3rh8S+heHxw
RV+HuWDaiqHvVkYwyXkXi+1CWXuWdIMjep+GAy7FV6ulShmqZ3fOtS91pDLYPDaCaUzUOJe2GBBT
nm3aLSKOlGaoJle9uIXCOsBsPTU8FWn5kb6uicUQ+R0nTM1atzvXfPJxBEaCTJMQg9JNCzIf4GDd
LeO5qxIU8svsvy8HT3FkbON7SR6/13YqiUHjUr//kHHxtlGjg9xfMThCPdaqVPAqmyrxXUOo0xKp
wGa46I55Woj+E1d0TgE7f3pvoGCrVktmlW8hp3ajJbAmuGIOsLD3t/dqy9KH3YmpfyYghusReoib
L9gu5MixXGbzVZFQ8N+tckMiK/td7F0XjzunUDAECpqFuSYEWVyu3v7r+nT3NPVtcpRulu19APB0
u/+Y3Hi5b0djkXEHmyMHn4f/legrjZsGwaQZOp84YtmtLZK8SeBWeIvZV9GwjoXrUVu8cuOvU/B7
aD4aX56ktLioxBKYcHCITUqnVpgyawlNgwD/zQ9xhv8e3t64u9Jl1t/hfC08u7NrpaH1902e/Wq6
mUKXnaym+xoB7Dz1BGdXh3Y+yhMu+wnNSq0YIN01OwPxR/CCGU/G3wmAAinM9oFqiXCRDMWQFg9p
OmkaQMrI6bmTZBSBN3+MRchP7tg0Yx084kM2ak+iDUzvzBCNQuleOJ1DpSl4x2GQmmTSjGZRGzvy
UPJE7+FNgrp7FHkf8oV1pD4YH/blkY8+QoozvUEBIy/8Z7+jlxKmF1rMsM+RRGFRWMIssbN592uo
xduHWymjteU8oyNFdjxv32tTikses4sBS5Vc9uLLvOaBD+wMlbnEb0OxQBeHqkM6Cb5HamLcr9sR
xgdbsCqBLxxTeAozuFmvqAqVFXcce3Xu0Y/F7Qf3o/hEfkubqTrJxJGHfBZ4QF78PQOcfh16iUou
vvKNqRFCSU5p+g/daXIDyymO+bxIyP4igYIb3txQ3JUZ7+A13qin7HHFjJ0VBEugeV37z7cGI+Bl
goZGgtC4UOM7jQmXa0bLlFZKA2KHv06evuqJ11hb/2nvKvlszv4hUxBlN/6qwRQh2LlaxYvEPmog
2Cy1NymLytc6M9VT4wBMWoBzK+Kdm3IZWAc+rEiua55QXSMOKap+pyp9AYmPZkthNhCbm8vwOXVK
URR/pKSyVf0trp2DdyYfw7TT7CQlse+9kSc/jIXdSYXG00vmmPr2wNjr7l4O1OSW1AnjTiN6JnzB
dYIBKWJs+wQ5Ciw+jH8Ga+Ijm/2fTc6vKmU/m9kUERjAfjJFBZ5sp6EV3ixjNZOqshKmxuLbUYv+
3NCAmVQDYYHC4goL4Dy9huB+9AZJ6aC2baR+iSDcrqEvDUhACe4CX0PSdipCKovcCBW59ZF7YX9e
bJkdjGOkVHinT7S83UirwTGUSHlhk/XTlS8HXG4SFfWVQtU3wU1caznLdIGruZ314WVMiJ8t9EML
dYZfqeJWRBQU5ftVAscbIzcRrIuiqinqRHek9mZCE+q2Nw0OT+6lvytNJ1PvAzn9fYIVL8Jy8Bkl
ROdpFVxMOHjbWbSOAPoIF0Ylgwf01qfc7hfV/eRMwdtBNhuvSnt3XCxRhQWth4PXy4Xity5hAOo/
zN7LphjaoSwX0AvNtyjM/kyKzRGmLuo9ZNBJAs0/0wnid+d83HsIggiVB/7vnhq8RpLJLBXp+vdv
tKextxpvz8cI0szfqxdfosqqBRhudFvw0Jsjox8ZUFgmlAYlvuRklnv/ounZGH3XNW67X4voqBZu
4005l5I6hSE55QxFpaZxknJlsJb4U8dVBnDKfr/9Hw3+GTtFlCHlpfGq0kuw14vjPdEfvWpIMZo0
89c0AqiMldDMA28WZbGvdotnfqiI1peQIIdolZFv65VC4mHNLlLLNR36IsoEZEaRzEQ+u4ZCQe39
/T9EzfNU2dlqX7ZlDNirGstZvydg8nPsLL3ngFZt7ENpZJFLI68S1pCZNqEBELKQhkuUynC3tSpn
uOE5uAlU/c8xYdHrYpQbTcgPq4Np+nuaWxGCy3KOYY150+Owsv3fYDXIuVDG5QEBrvYqIiVVNtZ5
OZUONCVKBmBieI+xjrshjr5Hp6FlckrY08NVPEyqZcl/Nwd1b11f7JNgvkVDpdQ3egdGnEDi6W4+
3prMdJsIYBsE+ytBLFrDDhAP9nohmpv53in0/Y6HcyRq3c2Xv63OKsz8SqqgpqPFWnyTVeGKdix5
FbUTYOzT50CN9mlCq0fhlWIz0Xd1SxAXHTKMsZMFedOTlcoQR45KsIxR6z3D2F7nSxlVz3KrhTAE
fUKCs4Wkvg8var84cFAd/d8uG+voMThscCCD2G8O4YH+Grm6XkMzS1NEH8r7zQFEeXUYoC2sqKiJ
GabtiYsFW4zGUFPvgHrpmcln1wrSN+pSRw1xipCLdL2R0zNCn91kwZYRO97U2UH0ewcM3kjJiwQ2
5f9SV6es20aTzwmYKQM9/cQx2fmOiTo2DzyJjnZZGL1+ioj9Y4URMA7+awgFKVazd74tbHmdl1/8
xG1hrcbjoQi50pfeBeQ3ezbgd5N5QwYMpN25+IQaqSg66Q6IJLJTEnwBXWZMMrWPxSsI4oaUshmR
dA//FbWmfmWUIzgy1NGzuxnD7FA0vV5Zo4Z7Y7QtwQtZdjcZtI4B5xGWGdEtWg7Fc4lbp4bfeK6c
yeX3b3P0sI7vjAVPuWW85xmxJxCEf07fSwu0nrA9EpqWaDYsY1cohbkzMkJf7VVRF5xJNAZV+77g
kFHgbeA9AMjwiL7s0JnlUOt0gq0a4RBiJDkbp4tRqGS5HSTp0bWgOgw4h5OSIrsRqMUTVA9V8s/3
irpe2plN0wz2WLLBfObGe7DvISkHod1Su+4Pn/0HXma9CNosA7RtAuY81gkGMa66KPa/YgsUi8oq
ictfxMuqWKfLUaseg7nvmDC7XLt5RMeYzqgnYZL2nlY4+L3bZN3TzFLElbzoEY/cpSJbUgzURdFo
0poQiZbpOWArl/69Q86SpgxVJ1nZ2U1PbnRt/vVQjwEoBz1UOx4XZTmgWPMySxNYRtccqlh+tqPu
VFKN6D2LhXnIy+OlpNKsnXrftSMVDYLDW3/s37CizlDkiiPnjzCOWldLaWI/z1bsp/4Bguj+nsz1
wQiUfDUQ++aXEz7v1I5cVFFfP1ZT8rJYCbBo7okKj6UK+rhVMYp9Fe6nM6rkXxn7XWcXcEngfFQZ
JbR1pcDcdYWX4zYNOO3SSl4P5+DB4mT0YsO17cc31UXDk/d1mz1SWrfQBBz8O1nN+Ol0aBApOqE0
WLEXa6776vaVOPvt+Dgd7LS/EhOV8TbVqodMBTCXIXyi95gYa+E/MfTvPMvsbR7TGT6eGAbK47hU
KWNrzOTcZshhvPgarpVxY62zIi84FfVR2IMpPCpSuQGHXXjQdoAYkRWknpPev+D+0bIayS8g6Brt
KrxHv/woD/e4TWMP2h9ZBG4LZ9ZbY4F//4wDDUmIBQ9F4a9kIv1sfHinLE2E7gETDj5AzTsn56tG
xSLFxLqOuulAPC7vQtnHvU/Ecwg2kCC4czZgZQ8Xwq/rm3RY7DMiqy3n/IwhCY8xckn6tRo/m4Z/
x2PZXqkzO9Icko8ZkVa2YjxFF/FsLnlfho1IcgayASHE68rALkghT+VuO/ud9P9MDJ+fnUB9lxju
SSZ7gU8Ohz/2CC4RdEuCWL0kjchp1CNjaP0ZI67LufrBjC8d/1ZKZ4AY77b4vQ+nTtSwX7/YAn3P
MLNjEGbeONs0tcx3w7erdcTyvu9xIeP2DkFC8zEhkhKsEiyiX9huVmBIKb8Ufz5dvCZ/1HzGmGQV
DjLZ4w01h9CxyofBAmM70bHToFlsrevsinmQyDIj43Kd2iQcvgkVxWgFzTTE0pIw5N6bmFvc7Vn8
GN63vgE2gEJEFUp2KQmmbUNUtYGpkWcziHX/ZsFwOfdKmw/eQEoYSqp3NfCXh4SF3rQXrz34NDM3
y7ZD2uI3HZUHbQXFV8g7kMaqiwzZhP6VIB8PnXNZZVhO+/f0Z4IwIHq/SruX1UW0KIv6M/rGalEF
B8qtLFe/96dxnePv//PxybJJP7wdecXlO3mIksdIw+je/gv+SteISotRgRzl3dPWIqDiJihZE0rI
GRJ+U0zS3mJQtWUbF8OjkG3TZRpgm+uU2LkuSwXG7YlSRSXszW4QpOkYQG69+qCJzC9msdNJVzKJ
pSwVycZ12q/dEkYMqpjaHzKDOOOfRybgwYannhAaClcwAA2oXSbnZkzop/g/WRUcDA2tbiI7fthu
KpZZbpyKXkIwcXiLpsRjs4zzpafBHhIw1g3ZZFeF3EBcUvrMw/NiXnPEpFWnjIgx1SK5YmGmWB6R
t0hI8pTJ4/1Dy/WxdSBx3jGKL8AgBFfujdUmwbn6oURxMcd+VzTfEP6WejdUgcdZ30siMNiszqKJ
twUJan9xMRiZu3KvRYX88QLnxmrWlnGJOmssfdnpPNuEIr1W+O2hPhhcqP8AvAKkFqUoW6NPyvfk
OH2dQ6Mz6ki1OjoWZNXcf4M7HhPA0hfiH/CJ2eeicRKoZLLtrp0WA1RfFD3IU533kRBdSjCOlIRm
rsJZKFPQKZSWNMHlcbGjNB9hYSINsH//RnZlFdtkxszsS33YXBSMRPCndO/kGqmwSs16Ro6x5aPQ
N7gOweeqolFi7cFvWzTvP0JynGLsLUof+9BiykqcQH+Hu52kdGFqTXhKMie9RP5tle6JgZ7xezAZ
SBg2YhnGMhP1GGtll9m+Nd+pRUwqGaIzuK1f9xAk2FRxlHKQ5oSFYq0mARNLHHJ+7jhdxxXhTBwq
KLhx2vZDn5CB3G6LN9Y533M84IM93U7RntclunysiU3M3JfleVhXzrw7kjU6UOltpIuncEweqFpx
Uoljghz7mvDmNwLnfyhdBNa97f8Vh/zQAAoLP/zpJ+41c1qTdXg552phHcMSatDCh7V0Avj6zQ3N
HGY3eFLWnX3cDIrxc5n2rtJQWTjWH3blS9iBTGvCK8NzsblM18RUE77QZtD6r3i3H5XJrU02a5Q1
NcC7rLFZmQZ6i2OXA7HMbhHixCBkgbyhagsTZJbBNVDbfvtSouVGRxsApYmrmX8o5Kc8Pt1S595H
PY2ogKtAKQwT1C62j0OoCJf7tDUnqD0Vt05fL9Gy/vjY6LRJzkgreuO/lVDF/eVFlwdiDiDPBYrf
PyepZZ+WLwcvAfw4kYu8ve5bOSfau+HpcFMH0yienITXyRxx8hMlg1HoqB9qIr6OyFpNOAqTUIdJ
r5IMVKmrMsSl7VCX/trAMCpc/fdc0h6/fpnHimqIs9ZO2s+bXSXmnV8ilnLgHAA8nUyS4MXv7rpK
6r6OyDQZRJfIjB/xPtzB8Qb2FtOZbnMstjBBOI65Hc88qGW/vt3seCuMhPXubli0p+fOqvlzpZZy
J+LdS/AosclL5R8zxGmnOsyAGCILZq0GhCTue6hqPD7RTsmwzRZ7vNqsoHNV4FZmjRrIPhoLCME2
6D0bhQbfRbQa1w+PkILEcEflcvK44dUNnbJOqnbMp9yRGj+JtWcHyEw48Y/FwqKmzD4LWsKfLwZg
33E3DlfsIe1zGIXArObJCAIoDfW3pg9nLxsK9t/nqne8znNfJUTSMoeZUPom/tyCTxHb67Potnn4
TW3Wv7huKc6ZCCrdUKjnCajIZYikyLxTX1HRzAiNKTIOXV2jjjDwiwESPmcq35m6G9pCyxoU9zwP
abpeT4PZuZQmyPLmzIPSapinwns6KSM6AKgibvIU2XNMod6CFqFa6uha1rls1F9lP6uack0itvS9
8Cxs8PjZUJ1W/Z7UhNLccvFAI/socnQnqAnbWAgsPmfrWZvigCj43mr1RDGvj9Nv067uxLwacZjo
j4048RB/Admp045FF8sc31KMvE2AwbyWpn/tSrc4IbYcleDGRlek6G849tjMOrJFmt3SABVkQPZz
OqFou+cIUqTuqR3G0BaYeZUx9xQPV9GJXToSfJzJBe1XV/oiH7H9/Fxk3Nxlvn9TkgPj1eT2Ychv
Lr/kjr3Z/SJE5u9IpxVpKBolL4WW4t8ah67Ix4bOVSZMpM9IPUeDr9HaqjZW11fzNz/wTIbjZYXP
ew9OUjBON4Fcy42/rq024I53VYYH7g5w+NZTBcjxTrM1bZDiiQ/cPp9Q1FwEujz3EmEf8fQdugBW
RlrQQzlCbW045MONHi6WrI2ZejHDq2oOQNLBfK0ZR5/piZajSGnK9oQd7FIkIsQaUjfDg4OWLMjk
XfsXpdFTQVFlgNO4ddWhpyZcuCO3IMiT2x7ujLi78tjR6SsvLbcPpgwtt7xljpjZnS5/n10hJ6ns
qkR0dHG6yuq0XOJzMrxyIC+Fr1Tf8xy3k7Fe4gSqtUb43OVqpdhDLFoKWj9r1sDzNy/gKfU/8TIT
OexWVy5wGBUid5p/iBVb/n72Z9NMHB+fA2z7nJySDoyO8LyRb7b9NT/1xDm2ELHvCJgzMS3a3LRS
CthJa71OC8Z99rDgmWAayb8SQRt3CsCGyo1qCdGkNpxBEC8HoU2Dsko01LBwH0xGDCAyscSI5HOy
Mp8R4jMtlGfhmesw58BY1o6IdJmcGr2ampypfsj8H3W4qTonRh9fxluG9yuM5G9uD/a7bZ23E/Eo
7rZ3Le2LISKZjnOBfM72/5/asaVZtgU3wQ5FDzVNQbp0WH0Yr/TgjqLL1Z60TKoY+M9Iab8kQpb1
XWFeVXMCXLO20QlZSa4sEfX8SWC8BlODWpDzX/85xyK1SvonepqOX1nxRuRxq2c4HSQUzjH5gyhi
sn1DYZkP2tBSgf6Ixu8HFhAyWXELr/4dDUQPqrtUlYamDvTMYfrt73CCa/rkAfF/C2WIcpSOzVtC
PGVQfXLm02iSyrabPqwdoPsfGjYRIDVjpAEjl3R2mAf8tm1sHLFLG8r4cwuUM3xvzZ+tuDBFUETe
86jRkFlqIgv7vfjlNqvpBR7d3C2dtErdDNGDGr5v5Ij86Eo2VvWwvgIquLMuv8N/DF3Z5DQTIT16
9AwadxWbCr8HFDgMHrPIW0EzlkozAnMRO1jmYmPnlubMiFN2vDrW53pQvDahIOCAhd3GM+lE6fee
TsPEIhc26nGeIATEb2eOX6tcmW8VxffVxgmZ11UmtUNZM38/a7567UXhhtOIOivQ1XfxPNTMQu/j
rtfpLg+iba5Q3nGVac676HDlrDDw/l2aSlpcK13TWAVsyLfJ27534aGoD2khC19CycdimCjL6tsr
7yRG1sJC3eeBIBYDz3GGVfN0sifk8MLb1qooqFJrZ/aizTYQuL3hdt4DOx2YWpMQFpX1ZEogcEHa
jn+8Hoodzt0fvVAw5DTf20ft5IvE4ovH+bqC9XLL6xJkYRpijZ3NY+RJKCDlTAtgLMxjLwofLPwt
FHmQ2zY7PVlhyFuW4SRAZEHjFtI7a5WLwf/5Kpd6TJfW4j6+rsciBu3OSnzoR0TvbUYLNlnnYzJz
wEQlgY+nfcfQ0R7TZof+3B1uf0npkjwIC2I/DNV3/3CPM4Zs8ZCk4I3c/ihtAiknNzvtY6r61e/7
kZWkkgw5cI7M0bENpufGt6TzwpM2kmHhHR8u5RTySNEziv/aMTllHro3CKQIBIbKlP/N3LeHOTeK
D5t0tMnkP2H/nZAcyqPRKKfeOHN2FAIYUDBkZjml4EOU6rkhHC9mK11zgFCwbN3YZ69ddndFQoUq
rLJi3HFHc9mX2aVVmkmC/4gLWSMq7VeIGXCrYcLqFgckHEnEUV51ujTqw78NI+717Rtu9qIlgCWn
/xdrT3QZPW2IaEg9v52E6+V7V8AE+9gTNbjFwZ3Um8vOKO2yNcklxsooCi3LOE4KiC/FeZDiY/AR
Cm7UMxQw6kjbzHRrCkzmM3z8njHE/O8OXYPneqoULmmv7/PoBsYXRaY8cq/QAPXSMuOafG+n3dO9
aSrFIuQjhADWMXI1DfBnsIPBWjAn5i3OVW7Tu1x8cGm6Q2g4muF8RNS2Xu5UX/mSj5xo5keUPmwb
Wcsd/1842Aym9a+8Dgf0/UNA6712TEy6JFt059NnLExJdJXQ4EnkH2kPUmVU1d/WZXQmF4+oxiy/
+mY3mKicu9cxOgt0/+4fDpHC4uSeSNIoc1HfAIZAz2EXrb4lAQa0+/TPcUGWbKDJIgkuKxbx5HYg
yuhyzcaibX6sizv95f3vcYMPbktsr7lqNVLOydP/PautUAmF0y7vubmTLBz4+CKhDSV1N548Jme3
0tmnnf3ugS6krQcR0AL8ygaSiqjbP9UEdg9qhm7T21MraQ6dDJQ6k1Ggph9lEP2MmM6IeZ638TXz
Aj4LE4j+kNPepPVbYzrhumM7Gy6RjMOKBnNahenMNtZw/Cirh+jVVDY/8S4wZrpwdwQBMZ7KrFZt
n6LsIEsosY66u4Qgs6SXsjlcC4Fot366ucPPo1nan+QU8Uik6HGZFcw/Q1Bfrn6pktqb6L6kgR5i
Mn02Ccr01xdN3t1XSi+f8u5oj34DIQFVCukZmAGmeAs1qahJj4ZRfmvOA1D2ogSsR8IExHS8X34z
hgExr3jKpE1T0BrT052l4e2B7HbKHqTku414eis/HABLOyX0sINCyOLqUx++7zoQSQENjIs/Cyho
6hrrgrJLYkMgWN7/r3RFB1C7ZWXI6hXUlafgLKT3WQE0LA5nogQKVeYETaE4qYoK+XC5trJdNLxp
ShybiDyjYTbiyhWA9IkEkannFoUO6l6G3hyTsgWV6EhaAaIlhCPqBIS1KPxvb3PSMmNbxQnoem+c
ZQ9MTC97I/MPqagpo1B/ww8NwzYil4OlwqhWaThba25E163PwHLfHfanLRZWQQ6yNS14ATUxBWsr
YfLquz20opRfdnhNng1w313k5VmkPb/QIFeiBir7Pffk/DSDLYR/L4D3BMmeOAUqAVpc+CKDEgv2
UfRCKh55Ygx2wejGz0sDwGmkikahhXWAZHKIvHrNSjlvH5kVaGEzreki6JmJ26L/TRuZHQswTqYC
MsYPu9JUKsmYyeNts6bEiytKGOqjfsoytcTKL1Pvf5/C6ujP7/naCvpl+HkSLlPzP5OwNJEc3sjj
hu5Yp+/lMiE2rIUpP/XG0QqEAMdrZeVKU2ao8ElzUHE6rOWeLZwvjtWMSADtfCiw9oRhnRxSe3FP
qPyoVEJlcXNv5ulrB3QPQ4Cxlf3JoOtJXcEi4QqP8QlaI4Q3QrwTy8tQ1B9SAHBAMhUDDpI7/OdD
ISsVMvLPAXVtfG95OlXDXDw3404sDbH2ErF6uLelJCb+x9BMdXW4SlJtgrSEn5M3jDahs7spxGVD
6MHqjWy8BcVRdAhemrbhUxjZAesSjbjY2jK6e1AhuROzChP1nAgaqQODyGFkllg8oc/RYftjCcAD
PvMnIQa2J7ySmulRI6Ii1bNlHF1v9lEfoi7Z3bzsBIeAIz0No1AmOYlMyEvs4LCr5gKfjAmQ9cpW
S2ZBGYwlKWH+TTeXsb/9xgUqbplYSdXFGWc7JUmNqtZWaQs2akHFdvOALDdZCuWTLDR3oOyjoLb6
LuYMKNSWdWtih364f5wtFE9VRvF7htCF69hEygfe+giWrz7ZIMsSG82bFaoR8ntmtfAEOnsfV7+3
0T0LJj2jIDXtc5jkhlqm+3VtNz2hW0UdXSk9QBrh+5ysB4AgkTHktYdNBNIOHzV16V3ZYyJpdkmP
zhNhzaZAzv2G33fZAVJfnNX0h7hQW2Z53XOEdnwKfanzhCU+LxgpquaIZyt6DNRf4tmxfxnyzSlE
D9NQ+ImNVJZmg2Udz9136XiqiEwKIQwSrhsM5bN4lebE7lUdzkiZYg2aKsvMhd7fq8QlbJFpkpg/
yE+mb/yE6wLAeGov46LEEpWYzr2u9mIKruTWcVbr5g7/3Ypwnyg78S36CkP0FNUtz4yosevK0oLU
tXJd0LrXeMjVmrRi5dfuL7AdjWyUDlHztACjyqMLuWgTjrHMnPLxWqtOPXsP7FAE0287ZlzHdOy1
zuMk9GE3hfEGTHmCquFTkr2mkl8RC0+3WU1NSgLsUYn2fs6FcJK/xdLiGwDEng7GfkB44CKvek0N
zrV7nfOQL9ECnywkiRucbRxKDrPkcGn6LwxxNYtVNpTWI4u3lcr+wZ/P/ln3CqQhRR3ANv0/JZ+c
f9ef7/9wJUlKRtVfd9jUy3Cv09t0lyPjgs939jzvB+USIaaeB64T78B7Ao2b5ekmYmfFoTmcN57m
+ZkYEgAZUNGuLJRj88k+KUb5rGnUf7UBouyLP5f0AMGx555i4z+G6HJ5BoklMsLHKDRIskuQA1kj
HyuSj2OUsfghnbOnGZzEabV+EuVVhPn/hQowR1kgv7iTFz9sC6GK2U8ygjgYlh80kCr/Iod6UdSG
uoZEPbFn1mbmnn6gvhdfcCj8kkG+U8D0fW/RTmheRVBhYmbT04dUjzjet5ifd/0iWqRn7+wxr3AA
+d3QVuaru+rx8Vw0xbdnOCZCcsUwjHsV7Y0sC+iZ3M6SCBmZJt2FM8rP5GOMkMZ08N89iZiUS0Yd
1i5bjC+3Pmisw2kci4HdyL4VuVRAmLQV1yD5HL9rLkMlsTD9LK6X2WqL5i1KhPCPbBcc74Zx+C+7
CSO2rq9qiML8gGIag2EuLXBBHaje0bKlJtLouoMeLNlwsSZB/f5sboPzs1F8X20jqpDoSktWzMer
NbBk6Bus5stgFx5L0VZXbrFGe1djVS/T1SGisksSo1tEC6v/2qECozBdnwjtCjcgOCakb1A6Yikw
XR7JSb04yQSkVE/9FNIhF3Xjjl0O3p519zuAQlfjswEXePJTW3VYhbvXlikTRXttQUsfBYoamPP6
mFPX9hsC0i5tGggJ9k9Cta4xca7kJD+AiRQgIeswS3iPHzxTh+5MbxM92ou60ALLe8MzMH6L08Zm
srvakXVLJBfuTCKGSfF078GQC7ZlaRDk1x2uRhURAmyMBZPzsbfgqZOtKYDBHUq0mx71Yy0PThCS
rZbnSLy5ljRoXiDykrNTW0koPKEYiHGKLAHffUcaZ6HJSajMwHsq03E/gncDN3mEi5Zdhsi2swti
ZrQqOhAF3CeEAOXElZoZQDtqx82a3tndsxL7IqLfa5ugtQ5b8VYCXHDOrd003MReXTj5FcXaCnKC
82GWJVDBNEXzUbqd2NCnE2+i+Z1Ruf3fSvimXzUEq2MM5Fd0htV61oSjr1J89wfigUg3wlepK8f3
ltux57TgOBvXxYjgcVNIZONTVUZUAlBZBKOunuJmEOmv36Q6bhepJ0DymZOS/kNwv9gDcRH15dT8
n201OzGk2q5W5kktv8c/aGcc5NWbYFX/nHHlYiViaZfkaDevhNDMmSSkWI+XbR0D7yYUaMP2OXzT
ns9enUjfAJwYRNZ/fSaPLwTRZW2m0IIDUjJSi3HDzermF5jK12OMXDJiaXFfs0O//CWWRKoWsmoG
03l4jDlrTPFZR+yErMIrNwMOh1cBpslLYlx2XDfofqFKHSgwJ3YaZHE8OlisNfCnPw1/2fT+tHi3
bc9kWOtFea6UqP8PsIFqI9SHKJD0GdjI82JMFK6kl2txkFqg4GM/QWH1oOu2BYQ8gOiAh9mEcdot
h+dvFq0m9WI6hmWljrfVOwlfkvQGLuX1vMUM2MDiJmxq1AcgqlRSXFeIFBckJktBW9/h0r8ghLaT
aO6rrCSQiF5IX+26i5c9kwpYfsz/AKS1mZWKduuo/IRl1vhWljXyCTMpaajJVrGYm+/Ew8GfzfHG
XBqjJqq6wU0NhtotaBN+kjllYsg88VEOWBWLkCDe/8EmW/xZCPxHwbGkKoxYph0+zXezK9tcpSyI
0XkO78zJzCkaML4sLtsa1Biy7KyerOgnp+u2hO8R04s3sPfXsEZiBSzF6Q0sybd84s9ahKkvNWCB
sQ6umEiRhbVWoUdNjBGRMHkOIrgv/19ohBhVMuauDh2jIjuNYHAJ7FnFkl0k3XK/3nh+YjDTIm3X
SZR6NGWoup9M/DXp6quzWQ4WWNnW5tPwH8exaXle3gYd7mqXDD93z9AA+CJRXZsyEBs2J0G3ISyX
McbwZ4UetW4+YwkqP811zJBJy8Bj08t/AM2P7FkEpaljk3tBGq1FCAA0kIVsxsAz/FFhpZio1lFJ
iVRiQHtQ1tHVqhCCSpJ+b3NwCH4rcwLWIWJazOdBMD7Bh7yFsxoej06mTfcWtXqP/g6tlC86PW3e
OrXjsdAkMm+LCSKKBs4G9kgI0wQwxCiWl4Njg9diZW3vQh+GHX3WzsaivK8gmmCqHimQtdIGE28a
cZjbboukwhB30RTxZ8EcHRukUDsXTpzE6buvs25WhTcaVLb953wBg+aeB/4Rt/JaJY0iUabR3akG
a6d3VBKztDezyhDIOUm+nXD+RXyiBPFwvNpNawNBAjPPhxZyaX8rbve4BCFMMLYKPM2KUHIC6Ffa
KpUwCwzty7A2fxbfPFjKtTmvP+4QV9IIlmvUzbQq/qJJ7FjxwAbBo0MUv45/oibrHyxofdMo5wE7
QXtbpbBSp+iFuGw1o3KFty4mjBfAfN2BWJrgcNXYLWB2vSuTP282liwkIbCZv/B67wmwowthJz8p
tpOeuaGKcNX3WBADb/l/pJ3hqU6qIcriNQzLB/BaOJB7KtbH4SyLcCfXHhOdtB7Bcg7hNGTXXp1C
DKbdtsyXDiUANBeNggtXVGPozO4A8G7lRlkbKRueXFRZAJciuvAtoQjlhpVlM3Fd5fu+gvIrZPxm
htCr1s/tR2Uhqs3R9hiElOeHEdznG5qHHSynpNDPapyEVaiZO6h3DhA3rnatAn7abAqCWncwE3I5
nNzlFvaQeJFDfTenE8/uv3l7CEfDuwydCoAeTbZPXYmiX/XeAYAevTSsSc2B9sBFb3vJNRRR3kH9
UzyUGB2cFp79O5qJ6hu2wt/0G4MgK0o8VVtEMqfOL7k/iRit3pVbfGqJLEXwGPqUHnex8IbW9IPh
zfCVhCik2sGE5eXCge2qJgeqpjTVLC0GueZf0zAnYvv+5V6aMiMb6yXNGohKhqxIvKisBSGjZqgd
Io8MIcwyyseUShj3+KNLEGjJkGtxELAwo47a4xdlixn6UK3cW3gnvYTb5Kg4WKE7gjK/In8+x+ui
vpeSoGu9v1cGhYbbIgpnmbn1M+e6polUozdzztrk4/5NyNbsrif7BbQypE/yXF2mB/6nNPj73uj3
i4l1RPsQrmQN4QCs380NN0CrhyHp8e491IBm9U02NyQew5a7fDs7jVIjMEUqDh0XudYVaw/mpInx
m+Pz6m8aR/Rs8QP5ODkLSxnzS4nsabQkFSYoYoIp85Grbdg6vgJVfkBkGhP9Uq6vsYhAQvhjkooi
Bu1Duf8uCQGtpxkad4cEcKrbyCp2aA1ChKIrjN8hVcypXboJGIkMYJElwtss8yzH6mGA3GNGITzD
b6cZOtmIa21TewtK6mkuHW1Zr3sdW1Pas9FPG+QCpFDgyPANC4FRuKpQFzPCVCXsu1gj2q7KdsM3
VRC5/8A/kUpCDqq7Z4fCZV8o0Muv7BlbBqXQFC9YTyV9b7nhBdpZXUAZRo7zOnnfMWkL8IuGuruZ
uBrJnybDlvxPeIA5NCP2aR1RLiGx3a6h3/ExlAkGlaAG14rFBUSLLqn8C7S1ZjXp7nBsqlswMcj9
7qQBemEnCMSXniMs7vyEwDB86ScjJY/okEDT0WlZ9KpR+lKn53ZF4G+/n98U5T02tNLdqCk663mP
SOloBnTx5+1JEucnenIwIRl/SFLN01PzzbpE8MOvtbU/1CCgnZu3XajvDh7ilDF2EgxA0uZ6Q2OM
tmHjfviO9zG2UCd5bfZEeKoTmqnU8cZXP9sO5egA9tBCC8oMXr5iyQEYHbiL8ImhylJu+TbKtvnM
Spi4u0PsjSaI3htri4AxmD7rwjn6ITJut7aoA92sPONN9I7ejAOjlT+53+AJXqHQmcyO4UGy/W+J
g89zHz4Sv7De8NcOT1jiIho/Ed5AJ16Q0+nF6P1sOy4bvNrpf30AWh7qH5V5IeNnXPZEIxoW/EE2
10BuDVQfmo+aojRLHWVwrDYsaYzCjPP+6wSuAxgD6RoL+tN6Xy1pX3yw35W1J1NZm7mTv37TjYN6
GxRsa4MDV+yUosLrNiEQl9UaZGb1ets2ipjV820ngWlX+EXJUXF2gw38OEKT29uvL8TSj1CicxIZ
iPedYlDx5TgMC2VosPL+Ij/TwvvT9Fk8ieBVpQeDxALI/CeFpe9ztNdt8wxJjonfiTMVqSIAtRU8
blDUkKzf7u4EpW3rdSJJ4ZZy7ms9ZkQxQjnDOMfB0kWQugkiPGU9VpeSdo+1isfnrnv4xERLueQW
00l6ArQaro0mBqEwSKjCdEzM2jQDpgSDJ71o2tiN1rBO9ZrL9L+b10DkWO7mITvVXh1p7HgSiXZa
j66v5QHIV7hKclYZhE6xSicDX2bZkzxSvMsCeYgs2AZVTD8SI/BiElM7b8+k9HTh3Su6dQvXqNMq
Gs8AcapzkeAyE9xc0MvA0pLWGQS3isZi8Gj5Y+BynmlnV4OvOE7n9v6L4cwnOHacPShQIcwLPAGH
sI9MJZhzuzPsOuNJIXPb3k6Ay1CmeZl+FN+8P8oUBNaSqwrzgKyoMfIsD3tWu6qim9rR5m6Jo5ql
7zdEVpYknckHJBTk/EFTbJudVIwndcpFxSOOsYMF1UVdTlFeM/SWRUi4+hzVz1KRp/b7yBMiKKSJ
KEoNskpylrAyAupViTEbIsMqAmwzhPcU4HQTVcA2V3ybal0n6ugrBHKvbRtVhFy75Bln9En3qd3u
PcvT6neehlhiO3pjLUbZr7jaejWp21ky0wIqF4lD2TdFw4nhA5P1V9kxUdhCEFAE61EG8PH+7GnE
bfSxWO+93FozxiNHgq4WemHoxEsUq1QiHRLwdPIHVFrxytHM4k6Z109zAblDQS5BlsZ1n20ivR7Q
4SRkFHGvg6t/Oih/SydE6dNo+HZNZVBQRbte3ttvGppSaczJFNgiH2TlqHX+aqTqhrtxXOdkn7qb
shhLJG9+17qddiu8Yh7NO+/LflgkK9uyYbGT8NlG1Gaz5wPCORApCJDqDkN2avDqqz1FRXipHs2W
EUdHAiMh5prcPp1vTNqfNugQ1gwimRy3bw8b9ReATvAd+WEBf0yrdbDZrIMWnY/tn5TO7oEEe2yp
ulylXP994cMUPGHL+M+5Yv62DoscEcSshfoy+9ZeguBvsmvqxp0izrwEiwDDiPcIKZG3YdMX7IwD
tn9bAhxbdtJpuSGuYDrn80t20xyNmBjXcNbBdCAIdi/nlLfn0hgZ3iSPPJcbtxQpfCvUrN+Rsmvp
U/jRJmg9OiYWblqjD/9jM7S81OnqqLPSnZCbxWhR1TotiMaaOJsQXhBjjvqn6ZY4qNoia67Jz52A
Afnqmz8t64hkZnXZFBFz5H2wT+vbiJJr7O7Vd3rhRj05/0LBD21yA5oKSEHMjGYRXltHoo39BZVW
wt3jyDUYmLtfAl6hYu9TF2ueDYJ+ARwWcKrrlIYH4EUa0iHIP5IAAUJREDha5Ez0ydyaPNrQUWek
3NWo1Pb6KXQ3a1AH7O3mvpOesRMs5+zSl3N3m8PZqqBPachGe1q5Az48Gh9R7bAqW28jc5OY4n8p
hIzhuJQdlgxO0BmOyw/eakmSzOVzSXDkMHKqfrvo77Lw6cvkjvkH2y53+9DE7bl98WMdSIgRlk7E
Dwr0KsGC9SmxEJMN6WP4q38K+VoNtUBawmoC8zkZyOxKdz11KCNgVqv4YCE5Es9NEusq31KdAy/O
OVn9RhFuk+Ger7X69hKBoBrp16YFvUuhDb3G+Jir6UK3f4GEbdWTQfGbWDgw8so0wlEB9zEWuJ0A
RgsTvrcvfdCSTajWNR8yeoOUWEEdvJ9XkEERQ1rde+hbLDNI+ToBloMiBpkXxdlyPsqoPqzR4rhp
MBmSA8j2vFe9ej6L0MJwp8nRoCJoj1SCgTLZNYBYusmBTesruhYk5/kIWxjC7WyVme7xTfZb1SCP
Hg6IWZp37X7BUM3d97dsMnZE5VXBcefWYC1d0FEZ2Yyc7NypYurg1AywZBn8iCPi8GOVx+nVqqfu
mQGOC/08A8OQiEWW/WIg/6DeX1tVwb61TCbVSXtocChzjNUDHIS2cHQF/OffbpMvuevQ+ddM8Z2M
X2w1VIV+pAs/e419eBXhnGGuQ6PcWeCKHXiUXn9oGbb0vmoIaFwP/+aFnMwy8OFpmtQfHngUu1Vg
QrW/eL6Kn/Oswp5CfOVKljaolUvik9+TawZknDMS3pD6ab8EqcaamnqYsQaZbQW7RNGJTlturiG8
AuAAorCQLm+ckzRSqkkmAs4K5ie6Abhxx977WWJe15AdLFywXBwpuL7de7Lh6UQRa1yjZxwOZlqc
IOv3xWgrMWyrk9lhRD1hS1rNLBzQVcaTQMtABVr/mMyWEP2Upm4JmZNWGVpOmHwgXXTVo/4j6Khu
jtGae+1m4pTz3wKiCK2kUahohJT7lhBO9Pqav1PGyjbUmtbGCK3dFj/yfjCvbWSVaeybmmoyYGYW
7kBDmdCpSCBFLZvFclu5qAGkS6XJ/s37/zBWzK1tHCUjiwtXwf3tsE8pb6oqOkazOI3QB9hUk/AX
s3CDH3vXXKYGxrJ5coNUUWtAg5mUbtJQ0RlNId4zCjtQU3YiskWORNWaFGcl59GLNmtChowZSIth
AHriATE84q7IF9vFmkSbiXxbQd6yCFhdYxMjtugX9QOsgabrsWI83lCZyWJowRhsshUVKuxeEjGX
tm6KirDlzyD7KhcfQa7T4FaGEunlJLscK1A+XSEPk/+YA1joeyI7KQblwHs5Jl1wCD0xaOlThUd0
h3aBpBKUEdfxMZWIK9t1+gmBVRcn9gxuwJsUyKuXaQwPabwaxao8TsdNixZlIX5SUNkwPBz7bgfU
KBc2WOMpa5KtNHdTS8+fvPxtCgnwvBttp8pBMkD2z5w/Z6bC+KEOkAkHYOY0v3VQbID01DheWKvq
p6OYjak+9b9hEV+lQwzUzVLHM0c16be2kfqTqcOnWsdlo1mHQEi/cqDOGvrNxRyxBY/fXnKd6PwE
iqBaKwIr3QIPOYVIPxc6LndBuDI0baro/QJn4zk8lDhtLpPaR1g1IuLjOU30i6QDeHyLfXUO2ssr
LSO33wK5tP2Kb5gFqZ0lJPzqeBjm0XQKNDiZ0bz+49AkGVdDRcLJjKaUDTmT7bYGZTfhgSCpm0GF
cA45ww1FG7T+xq2ElVZPc3U79BOoVe5QRN+hPUgrnW8WMm2oGqQ7ToPEk37KjsFT/5+Cvnpww2ta
l6KVzoQmCXkmCc1wrkIz3syeoJJxWmwzx7QXaWj1OTl6dr1IEdG/tb05zp5Su3A+80LkeXNIzwDo
Co9fCW8w0YRfVPJjr/Ftso02lzcedLR/nEHfCRwbjzeCbrm4MdiebeHAAfpXuyBP7X9RmuctR0qI
MP8fNyDhpwphcACFWLlBfXYHffLlHzDLCQM/+71W0DISLCuaCdaGQCeliTZuTFJXaFyP9pKL2p8l
b+9dV4nPol0QSLTZQf+VcKe/5/pUFLsMZMQTGq4IRUyi6XzAhSVjOqyEjNEdkU2RdjqCMJngIk3N
xrmuctF9gSq/qdk/Gp0v3kVTcev23FttB1j3qcHSbUwPToOC0A+nJ1NkgRXz0pQvCDu9crUzdATM
cs9qJYLhMxyQZCsHZ3BJjF1RmANjVjifE95mx6S9GY82ltMCnL7E2YwUK1RRgV0jGYO6JhgSnebR
fuJ5RQv23r+YpbR32HZeS8zEOOC++rP7n2m6BhYBZW6T56pOIFGQYs19nIWJK1JyvwuIAXBqCaKN
Y4AzuPr9+yk3ofXqHsk01tNg4wMhScmiDhvG74WYvvhrp3JUtpCIwAqoXhrFduBS/U8niov2nW8k
glmL9Nole4OlHlSWiqBMX8Oaqf1BfeAx8GZRKplMvwEqlJNGgvRFi4IYgLS/KI6LCQAFfoWsCYXW
hM9WaRa5r3kOrlYSuOmugl1V3xcMBDkiwUO+JGOxpACieOLUGs37wxLVku+xm+lOXdUs+Dtjwn+O
EFsXJe6hc1aucaARhu2XD7zseRhZ1tQRXUV03jTuZ9pJc6oksKHTcxYlhMZnFCHIHFEWBrcOm0WY
eP+ScpoSyWM1bqXXXbvjCDjKWSFC9vbhmA/hJXvA31zKhjurAWojTyUAg+nLeppXSo1ILsF1MJ+V
0evtm3UyPs11dchdhfhzR88cmJ0G4Nj3e/4DipzFVJAeRdu0aBFX1OWZwrDTc1ubuHQKqf3PIHXk
+KBRJTjBt1fMubHIXUdIPZtnf9xf4cSqzq7H6AQ5ilo4IvpkKRe9hTThvFWKf0OHpVbsx+k7Y9n1
hQxjlExjSf5U/MOlFVGutnL0WB9AAIN+h5nA95KaGuHJfTDhdkdKNASAkiW0InM9YIICHqvleJYE
0nO8tVKSHvE6evqxPPE951gk246aKzkWTXTAPAp7p5RomITCz6DOBYdxsuIAlWvlTEwx+hhoch+W
Fvp5QMm2b65Gg33/aXrNJLeRKbECM9Qdr8qpDXogWSAKJeXjff5BG8EQKvDqLAjAYRecJ0qR5hMs
VWvYZO7LIvKgmEeGz5GkMm8PtlC6dedbrfcYNhfdIzOry9lOaPfd7h6U+p/Cp3ygRuBL7ZFA6Ru2
lFVdQSWxPsoW7/7zaPNxSITJMj+HfgXhd32MJmu0Om3QUhmfNoeRtXWwtABXZ487RohvXZyTF6uQ
c4QVYs7kTRa90us1sRxqjsFD/HHRyzB77o54fY+v1fRTgt2ZvNV0pmkihC2txLoRYQdK1REhN4cV
QAGE+doZo6IWdztibwkPBbjvk2F+sVH+BqQCgKewekITBdCBWvx58LUolT7Glg3VzLtS94Zi+N7M
IgoQddVri0J4xma7gXrVDXCbT+qSa30n3OwKJl/FE1bxTsnhJeXA0yy19HoEEY2PCf75CiG0ce8p
0LtHUBxZWiwalzYrtc/tuhZVKCpoVtFyGHQFIPr+1GzxP/xJe0geBXzRSeruFEPwpRIRrlVZ5Whh
tprHDIVCkLan6Xt66SRkCB4aewyzXwlJbuvw01rouQygn7xIdFP5pAVB37kZaJAS0MXHzgnZg/dP
ey3+eXH4B1U2CpcZ3/EZY7gGQmwJIXzUo8xDR0MXGpFCVRAX7P9Jd+5xj+QnqGh+16L6q1o83naW
YN6qo+z+K1tENjPUGit7mVwIKUxvjCxUZWxAKFxEFEsYXEoZZIeiKTUv0DqX6WVf3YED4CR5nT2a
Sgsg/r/Zn23ts8L2z676GXS/gkledgvtEeb/wvW3wvNrnrYI6r/DrljuuGt/kYaqF4Ny33kz5/Q8
OpwbC/DJYxFbxR884YrIcwVaoclO60y5HJcHmKEOHOnW48d5gNcnHT2vzz0vDAq/YnHvJ36uA37J
+npnrTp935pmptGs+2PS7Ph1RX25/2noIAT0T7xro72EdZWCYdAw7GAmsyOb0KHN+3sLyRk4iABt
PrEJO8ARH24FWv/JittlAaf8HSXFP37BHPjZD+2VnHF9JcglbSUf7ACScJkcu8hGk6E1vK8qWraU
Z4QWMw6ODxfKEODD6qU3zTgnj74apcOZIsLg5AB60ONzLfqyNOQGW1M0vtd8Rlg4ozgD9g==
`pragma protect end_protected
