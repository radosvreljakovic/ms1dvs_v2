// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kHX2gNWiRwD62hN9dDQ3PIF8hrPBvSZOat++M1sPFwESxlRlDSFIuZbJKz/MhyGW
fdPbUyFSiKjDq6lKiXGG3xzZPN0sj18LNsWnfZRy5A2FYZetqfbRmR5R8MBaBRp6
sa8nC2GmxUmYCplTxCXb6OE1kjLJrcVPLuBuXKL+cco=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57056)
BZfMhWLd7N+p4+QFzdlHcmI2BrFD8ypsaCD20h81vv3KKMchQoivNa4spk2SK2u0
kEQw6sxhUe9rNgEfigcWknw6BSOeakkz1TlXeRY3MMk24EXS2+Yy3a5Hqmnp7bNP
wXgMZPu+L3IoefWZMr1Jnlufw2vlvmIDIab+94zfR0+H3w9lLbOcyPA06lE58pgx
FBChHqjLdLD1Yo0pTzsVhJh8LmMA3Ria69fWRyuhgDA6OCkEQAKqhZ7NOPFqH94+
0dq7e0VHUkDR64nEFjY0afJPPaL8TcC1QF4/J5i2t/cb53uz+BT87XRlJ09uw22h
DmSmShYQ2kCEYUNQAobTEq3AsOdOY6WFAkrrM8OJ1hguFyAKn6jzrYQZ3AVQ9pc5
X/Ce3csKijCoZhqPcImidCcl0nY/opIDuce65m+9w//j5NgV/+GBvlCSRsibkS3F
IukelZRblVclR7F/68lo/LHhf7o0dhSDLgFo9w+ZBdE85ODaChYeQTPiAgzedjU3
bxjtyDzEo1p8XWoGSO+xJ1U6JPkj+/yQhlHJEj+N/eej8pKCw/JqVNeGG6qW+M0T
xwpQqK0UVms1F3seatUzh2BPqCEWpiCgzPbgPyv9c2FseUJ2KVlASzcDApqvET8/
a5zXTmr4s0f7Soi1W11NsFj4g2J21/tzFzm/9EEpqjJt/n6PVw7nmfx2uYW8CT1C
U1absyFCgOgrlmlP0y3hkLqnmwhxjQBSEJQjTJaDQqWcI704hPw4wfuRUeIKgpCX
IozPWfPXqAOAp//5UTIqmQMxlkywfok4j9lglLlPAUFrxGpVLRANd2u8iUYg6IrZ
7y0kt/ihXnkhYh9sw4lbQ6u7n55DwhlZrFL+aNw4gPj66njzTMeh/0ePuu5EjiOh
1kxRZpkE9fjoZuO6/d5n2U33+MNQ+zVouMk18/rpHIomryNQzLmiDXOJWhNQWAx9
Ef1qM5YdMq3EJSGxsJc1Qygc54XzoD0FyShMDokhgcB+K1ikBnMDyybQ2PiKhJZi
GvYPdbfs6zU9SsJxZYMT8ZxjezpSmPtJ+8vC398/WWkAgtO4REU86SVQaNCgTgcc
Zk/t6x4QB8zll1n9UPxHvKKdqxZnJ+WXZpB8TG4zuNhzYz6xueqc9QsNtDX21Z5X
nWhfxkFJ4WWPU/PkaItZT351kCruxCN+BacEVq8CHzRSVk3DUUqCCrxKVAkBBjE9
emfYJTLt/V9Nkd1r9xx5SOu22NYJIenv9coR1gX+q5OTENNayhDSa3pqHrhJPKKr
Q/vwGxFmJc59yOKqXhHRlHVq9cY85kOpdkRSEut3uo8JBJHt+eda5oN5DiSYKK3p
dHFijwIwY0VBAi8fa0Y6SprLg1BCibEt60/GF2pnX8kJTiD+qwimUGp+Wn1BZccL
YQ/ihwSLmqMMc3fWm1tDL1dyL5wLItm/HZpU835CNIWXi3j0i7Mbov5FRQnKEYX5
JVhnKiDR4oeuJYrYtaUM4GKSgbuSHDZX67jaq42ToIxpPj2hRMVAQjPmwsqsu1RU
FCpc8kbZKnrSLf9Tk4s1/XjoPJ/jhN1LcgHxKSbE+NVMXh0lVsLUBBcTaraKzQB/
NqwhJuCaVQsp82r/inWHp2kiRIAFoeVlkVrs30ElmBA4uv4Y8D8srxf9qhRhAdNh
TsK7wjKSifPLUph8nDBYkNzX/TyAAzrlijWk3euL2jOK6ep1rrXoBsfcw9V7ruu5
bcqvidyl83+OSUrklUKYq+l/zRjkFce7OMzCd3F+xcJ/xaz3/oTA9hWGw9g+UsT5
FE56a5UMo5ZNSHlPWBFNGLzGIWKWfiQvAx0/lIGqX5j3Fuoi3IwF/KaRmVFgWUAv
imRnVbp6IGMOiyK9qU3vXOHTY3vn0+0PZXgaa407Sos+r/blFRBlBRlmn0ioehgS
1bnK+HN8GoNOkimMceOBH7TjRtJ7UYy3KZ6MDm2iS/1pvO0fZPktcbPcLipJK4e2
8FCSfbzeli8OmcAQmu16SyehVB/CAVh/Bs3A9c7nlAkhaSI7HRajili+I0Rvdehr
yH5HPBlYo+K/fzSfe1wwYxO8fArIKL2hZ25DTrD5WbL+uyXGnqfcvcwHXzVpvBLN
ObXGPm/H7uqNTO/ZMdf8IxBl/B0+L0INCqX666w7l4EBl0PfkqE/McOmjmxJ7pKc
/4urw7yHV4ZBH5n1+wdKjLbrNB1tzf/XmyRATieURNLN/YFHV1570Ji11D0gLJQh
6PdnGaZbXKnOiIibGQ5WlxFApUKxCfe0WHNFbzj8lQfw9ytC2MdHiwZ+ZbOcv7fQ
+v+CcxLVr9WlKThKNFKfXn3mnkt6RCUpUkSZL+Od5E4yAguJvDWeBpDJXzVxXiZN
cpwtZ2gv2/oUFfZDZxpsbhNXhUSLDAljK1Dt5vG0vlBZ1TRFhC9i9/sTpnsUrHub
pZepdwZEtD8ucUcj6n7zqNhodyo3qqIfZXuxWoju8XnqYjWy2IgE0kGqs/hDx9SO
C24MWoqO2qK4tyI/VSy7QrVuTK0T087rpW/DD2AtxWuru54fot2yJl6RRNa03GcX
xTs8jhWY1a80HRYlA+HohOKWhR8YpcsCjKiRbJAIWOtlsy2cZNId+QQ/FH0/hSEw
uqapEyUlYktMtQzGpbYomhbihXsS/WhnHEGBFEzgTDtQZsT4EU4Rtooe3UPUm1VH
fPz4WiD0+FR+kKdkeI2jtPuKke6F4PCwUq9Ueti3Y5CN5yG/rRA2Ku7A+n9VIPR9
Oz/3FF7X0paz/dgxDXKucR+lEJ3iEZVtMA0VXiNEujIypdYLXeg2F8fgzjo8BsdA
JsfBhVsJYR3Shx00Shx8DQybWj82c9hUuubf5k0LkQH9ZSGr9BmjqY54eduDMxKS
k38tKUMwbvb159S8hu7XblgM7jwGNbLrjsYhIT/kzR7QqOFpiINdl0F3DurKix1y
Gddmsi5cL9p2GzYwAhfdpSPSqzlBEid0+aeb/QMZbffggoDeEKiBnKT6Mn8UeoOx
uXvA3wTpVwMOXW0/JcgQ9q6GyJ/vEjy6WhmTNC70J6IqSsitPp9iwnjTZ6rGvRU1
GYxlzslhRskPzG2PV9ld/LtY8mgSMFikvj37zUkL18UIrGhWorv9pJA7dSDI27CJ
xAMKzAvRyQ3Sn9IJKt/3UbzrpuWhMBW2NYq6XjT41IaoU8yoPHJI1uWHApmXyk23
0Gdddgxk5sPwkhJgcO9AOrRHekbh06ljkIKZ1wj9pPKynl71720dakSpjhlB/1Wy
fNYUbDwvhny8+EwqJvZgFBE8psWTX68ZrBILfI1CBC7UeWLEStQdxj8xXBVTWfoo
t1JW75DG8/Y0LKRgwK748ZiVDx+VP3l1FKVaF/vqHXVUMfZqgmSe2XvV+hXK80kc
qKHouuYOcGRgieEaC/6qQFXtdbTYTfnhjNL7tsLpF80bTW/axUOXMNGfZC4MyBKd
pJyRG7qC+5E6Rsg94aCu1eI2h9/Fo4F5Ez9+neYofLo1Tx767d58Q9jepHfGPgGw
a5x8wrl4XCQQeHvu86GTurJA8rXGq/KyHY4kO6aTtRFy3E7/BjurYw5GY4gLUcHO
PjzlWYHFV7JrUaGndAwoMYDXav9LuL5BZZlDRVpwex7X87IZDLliPJBXVumbRRhP
PlE5wsjttfzSKhg0+3GC2nVCWbR4uyMVPBCkMYXtmbaI0bfAh0W7SoxZ4R6dDnke
i50N3kr5ZL+jqGMUbzV0gWSrspqD1KU3U9TezSIbFrKUkR/LW/MkE4sA4QJzv2ZI
pJsofaii2+Gp9mH512bMZ0yDZMxS/x66TUQEw61pUUqBTjjggl+Uc10Hg//Of1cm
Mo/vO02QkSp60KplVNsCMPa6FU4RwD4n+A8e2Q2m78Xxu3mbyWQDZNCc2K1JnQqR
5OC3Y5nFFQ/oXxoUOUvUl27NPLhfGlZifojx2mpC31fFpV2Uvn/lzBBOW6Rp229z
ycUUXH9KOqvtmy1aDWspwcut4AQssA1cM/mu+giNucbIsxB375cVm/mV4zWK3RCr
EMeEBL6Ko8K/Y7xDN5yDk8Bhpj/5ukCMV5QzhslsJiEDoqWrhhrJtxrj4gdxAdIo
BJ9UzYw+/pHFB3hR9LSi8hhwgHqpALPG9O05vV/YtVoDdGD0NcyylREzcPXErYox
FAHvDM0LwCmMGYuth4oFZx3k1Wm6EEiITonxBzW7Yx/n1TG1SAUWPrPrNFzhz4SY
jMc8NLoUFuAWWbFqPV0d+RVhnLKxOsZChFrsMeIfNnC+uS7hfTcb94YIaFmvzr1C
Jcelh527Yr4ma0t6sknmH1/35WBTNPuWPUMrOmbJtsfuuIfykxsrA8MqiYGPZQ43
2axz4huzn66clPnUPmT/a05XoGp0k6YTTS1sadVtAR2INTfXG/NEu9sjnSqpxl5C
wRseZIJFvD8c1qNhhAClE9f6lzviC6KlE35B3pJEzM45NYIuSBma6CttAfCxtWVR
AHWdzR+ThoVs+9oZp/lLADp5OYdksyZQMOhC0vyMt20VmQnyo5T/G0HSdr3kDFns
oIOoXizQW3NPl/qIU6803iHwXQq2qyxCJ0gnh7P6V77mI8AnF2acmj6oNxPWzt86
oBK0cyOrwo85OeHmhV6J4woOnReH/YMzmlYV32lpok3L9qCIPA3/N62fPMm0dU8U
Pl+glFyueMer9whQTSalgqVSMnnD0cDVXXHQTzrGJ5qlxucUN+pBbDZF+P16fHyM
u+jR1PenELr8ysG2WEZE00eZO9cfl2/GzEZbyXFIakY4xIs27tp0PlCtvk6HwG5w
8VjQuNHYRw3gQyE2Xd2zcrw4hWjjK2cA8zwJhc2iEV6ONSmqD+LNUZfEoeouLImI
oRvddBMiHp3zrEiLDUvWY+aPzkKAEh2KqVxcxvCpezKEtNHp3QzcaD7zjg1H30cE
NzEuIIm25tEOttjdBVJME6m9Myajm3FBllOhZ+uOiasyoFRisLa71jFmaJz4TCJW
nabVeZ1ZXulOBYGnqDEdRmxQcBFVObzs3V9YS7H/IEGJZxq4t0V7CeXNXZN1K8ia
xoippnqZ11cGQigrBhOcl1wfnfhIrTAjGvpmmjmZeCbfCx5Jxn7CllFLkQg6xTrQ
JGhhTk8M8LWzjcvmbK7ekcbvUkFxEPnH/TijmKIMgUXUPNbsblOP6inwJZb8U+lZ
TEjD7nUYWrWQWKNJ5lzYlGZYaKjGCYB2dYVuaHh9Vc+PxAqdEHch+SbAzx4ShRKC
Hy41WhDJHcRqP+PLDQxHRzSS+DNJOeaYhxs5Uch5+ag7mbsnzREXfqpvMGktNENG
u9CviS0FKjvrXqSyMaURSJUmT57f/KKrwtG9TTKEyMtCth1oGqEPLI67ZNcUpjkR
hoszv/aQEcebSoWjlB7LqUe1x9LTwtKWmCXIJ8ZVAmvkkffLU+FY1ReJK4FqG7YN
vMMOQScAEedLWeaf8K/uB1Sb/GuBdBzF1tfxs37ZaDbFFI7+qS1/c3wLJxvN36bt
gSVdPBynDP3dy9Qb2qnOlx+gyzVMZJup2j7zCBn6TLU56jVLw62+ylrNYzvNX5D1
7XleY4QONSdE3pZR/S3M9NkI4nx17gfE5hIw2w0q4WB3p7jZexaXuiEarRJpel4Y
cJCbXVBN8Uvmzf6er7O9W4Kl5QeeatsCT0bcgeReeV79oqAMX9sDvMMfL/mZlf6z
AXgLXjivzj7kgP4gbllmgZj4lh4+jsmypFUICaEyU5iMVDIT/vZ05/CZuuCbLuQM
4PmL8vuH4jqmS6DA/cFsLNQR5cvzzp+zyJb0T0sCdjOJgKUmVBng/KL9qwisVbE6
XYRA+pX/GXUtsShyREmZfIhNyWzNOVpZSpHrIVO8jKwVRFdBVSygiDYMGx4KalHg
XicTv7KgODCYShOftseFV449Lya6nIIiwUqiku5q1alq5cjAe09nP39tFwHih0Qo
VCt9A9QRP4MS4S9bI73HQ7jtutq0KcY2YycHrcnzxwxTz34bc1f7EpG00T2UnGSv
i0XyuS8qUi6JOMJQ2D/2kWjAoCCgad37N7DC9UyIbiuFGw+NdK1Ass4AF0q4ELlS
08/dWzMdnPaFkNjbGLzoRVNzTP+JKP6p8PsyUdwHB2zElWYIo1l/0sm7T5foO7hk
ckSUX6l0wnBxxJQAflhqWL8cOlxf+3aMdepAKRP1zsgESWhsxoSAwsKzhmEzx+Ba
B7nlQWTHNhe0q+4Pe2gyiUTv6IR+gDx5m9eV6VNiip+EJ+HUIcsXqdbuf9/APxRe
6I6XOCfwC14bJK5SpgfAEHhYU7thXKJKsp2f9EalX/TvhhM/auvjpYwQRRZ7XHxo
4u+czbT0pSAYvH08nIpe1uQ7erDPazXuw8JSbNdL8kiu4aass77SC3EdeN1X6cma
9ldcKEUbbiDWLEf9oZdpFybY0RaCqT0VNoWfMc6i/0kQCcfvy3UDLCwNCVK9gIV0
fVWnaK/1hGIFGB5R+fb2RHhdWxUDq7LHIjR5rsiysvs2OZUAtODT13hpoeTbF6KF
TKt09GjRzRZsJGZvi1OKDiElzob0vbA0XHREZ114H5RqXXJqsf0iyY43cL1uEKaT
Eo/3ticB/Ew6EdPQMAzQUVTVUqK6mAB7ZXvCYfOY6BnRKwT3K2wYLSpxCqedlome
Tb8q43R3w1mwF2ekHhjUNmx52b8q0YiXbVvmBZljSAegx0aJ1/dmcj5ZUiWURJzu
kHTntL/WXw01qdAjNnCayusfSWXk6CWY1/fLZbtXh1hdVefbFqsJp1ILTfKue/+R
+SoqHeabLV+kYIu0BRT2rdW9b1aWqVpOCmCJKTcOwmFcKTk1zB/BdKG4qmPPGFjC
c9GjA0qjlqpqYwR+dRl7kxlkRhgKNIsZyBKhzmJc3SQCquIbQImsa4je9nbqw4Rf
xlwgCjeItcY0is8jrWc3VnzFeWSewoz7tLzgxJXV2Q4wEbWkEGizDcqy/nP2dID1
QBBKwmem08uL2W5IIw/DlaLjEg3ldeH1/Gb2fDj8/tMNS2+3GX8mNB88TzZ2MFz4
uNS9nwBncZspLKGrFMxtscth+NRcVaH7Ms1U8Sstokee41yO8GNSSrDmH+DRgS1P
md1hKvBVSy2XVH/q2VtS8vikgcfbHXi7go2oyUVS021397XTPjhVSwl2G+lMr5Km
RmnCfeR85WdoyZtrUzgQJ6CEC+hM6aFc4EaNzKdwmBRv/4C8BsOwixVCFaSDt9Np
DZTrZ1QLMouxAf33h6Qap5tWFIyBRJjk3tng/CUg1fkFt7vlQ10uXJCAL3UgezdY
+FFXF5UJnU2iw8Td7EQ3L5YvLTfooP98GoQEEYypu+mah/Lluo/DKgv7ywjWNDB/
+hvn9dytOb2bSlHDHxxNCk+c8H5QI/pFcbfqgOHWeLw+0mzcXSSNRJPjucBrMvRu
v8Hux0K/UeYY6Ks5uNAvVnCn5W0QPYfL890ajll8dOp2cw6jvSJ7ff44lDbqtwzO
XVr1eUo+at05cA36OlUtJTRWBLyKZmehMXpKHteJejlj9yCrMv1tJz1wDxFkawS1
+NYRk/WrQ/Bk1BWjZuVRxNAH7wdkv3rzfUYA+1YwIiIi71wxV7dmI1KL3xoR4Q4X
FfU9oNEOXWg6fYNQP1L2K/jx+PuVXdl9nlwgkVj56R2NRmpwC6qbrqSU7mNz1t4f
Eb/x+sH0mXMQ4cnR15MwcrcaoBFDcqGfkJg9Wz4L/jHqOZ5wSV2nsPujYwHopA66
vzEDFOpuqpiSINEktMbuM/ncugLCc27lqoWMZNv11zmx0YUymxRJK1tZXF8GABXX
LSi49tDIVnTwfsxrfC9lnAHk9QVAU3k5cDNoFWW3YUdCmdQWlOyhEs6EMkvkPvmR
SZ4mn0oQ3SjowkcU0AWP+2JwearanY/SpDAb19jHGW9lVjS4rY/TG2/mI35pQFBF
Qpa2paGxhtX2U6qnPYthsj9WvTK/nlqcG1WI3vCk8Oxy3G0NY+W+5LuVKKMHMycv
2WQ4bxFWaL1wb20a2f0ueXyJfqEuotU594+V+ZXXMx9lTdPhY92BIRY/FQp7yxXX
m6BgojIU4jgFmHPnkgDacoQWm2yAYTnYgzc4mUHEqLcYSGGeI28DQxVxjBYKlAvV
vZsuBR1YF2idgLL1+KPK/boeLPSnJQvbUK6SB1eXFbE0EHQfje61PXhKjg/sozuT
rdkaw6dZyyZm1okiKsn0pC3nm+cO9nQet1KrgZMVGyEIJHZ1AnYn05TKTQUwwJA3
3vFYdk1m6lCiHdzMHj5Fyy1C+dMUdkPSziQPrHR7s+2iOM+Lsbb15m6HmvVl6O1N
gnwRw59tr7nbthR//+T5BjRhaX3KJ3Huu3PXU+ywslnlUWpKhbJpWkQXQd2mMrgW
/xYl26cA4YXQkhmwNnS1Vh4MyX7sWTOlvIhRKrLe/UDAoswtdXR5B5qDJGu+SKVw
8fO1BavGn7X3iG1GJF8eAkwnngufBx3gh3jd37c/RrsUCOccTl0Wz7w8cIw3wNgD
83cRg6X4ivqGNXhFWo8HkCx6JiqB2Z+vD/h+93vGTKeCrXmOBnQf5JRWYwOSIv+Z
vs2VIy8DJhvV51qOEMShCFnxtP4HqyLsvfoiJFFuSn45plC3p+PlznF3W7v/Y7uQ
r0kbIU8DN97GgRiW/CvAGpyFd5LiDny94HYGwWTrn/9FZ9HfgQcrtD8PH8zoT1+c
05m16ckCxNrj/nPRYsGb1cnW9yhy4sAfKbOn//WGi4K/ILEp9OUEx7HzpuBjfKp1
S8dG3D1W7tELQcX91MvUdEh7ndJnEYSK8EurKyEC4713k2kFmqSMvg0QEuUxYrCT
vpwl2B2o5E37tgQH76K+rSFZIZjQkXhM5Z+/w0eiTgtf1cVEx2GgiKbQwxLHCRDT
r4hpfWf6Mqnn7egSTFt1BjN3nFPVPA4Z5LhUH10DfH6lhihHm/crfzeo20ZyIIgP
Mh4YASqtZTkbde6z2WLgpBgO4xvT04hYxjiHFsdb2KG4rkNrg8gF19MWCZnJvU45
GodmcvCM2387P1JT8JEbl/fom6Bt/Ymi1TzNu4h0skrXugAn5WACrOYhLVQjOHSd
GygwNLGBVsKkm1SS049yJHtizTNMiPblix/SAUYgkEkEPCaW0laqb4RAMTyPnRpR
3bpEU4xAhoegb2xBTnVdxl9zjB5wZdNltiExXaUoIzYWF6jObzBsK4XZcHUXooU1
FUxxEBxijIYx87jogUqRDo4MI8l0klgbjZU5YlzkYSBTnPd/S2HtrLYN3XaIgVgs
soyEa8+vClEFV1g+dEdF1wfjrnbReU/VrxTyP9XL+BLgqPbEz05KG+FBTIjv8QPw
7796fG/ihjhJWNbzJ1ocsumerMlNHDp7JeJOej0d9ZZEwy9lPQnIWw6oK8NaSCHx
eGvjUFyvKbbYU7GGAiawE/8VQk3yTjIFEoL692D9I0wgTHw2YqkOH+vQrnjzAxlj
ZyBZe6hD3B208ggbvr+NJeDkprRvTMXFAZRg8ZksVN+/Oyf/HmfVc9ArAbRESAvM
mWFEw3hh+CVB00p/zmxaVPBB85XmMsUl0/AyykKs408iuMpx+9QCiXNqYLcG01EI
4F7Kefc20vxlwryol3NU4Cgz1r7K82d+Ywen1/HwVDslf4OXTSKYs2/5ohD73fWv
DDeeHKJ4PGX80IrJGocnNt7CnS75KEcTSTcI8ILOQYdBrMe15IZl5mESKHIlxjPy
nLVhaWvhU67k55mC30hjaq3W4/P9vKFqTcu0qo0JYW43/zF7yN19t1p2qSyg7mJX
zx5+GV+zA2nnCFM79VDHP5WWv2lAiSXR4HyR7BqFHWqWu5xSsKhL4bTmxlhAuOEY
AZp93OxiXx6xsm9hs5eiuAZCREF+nW4YbnTfr+/qvJGs256xkzD+xldDmALFlqKJ
0rlObmwOYrVkMTp2z9FL4nhbxhsTg9fD7NdHatGxklCluXK5JWDbuS3X3BY7Hu3b
LeFSpJR4S2fTZFW4LF6Vx/tZZAlsIKDfPJ589hfe9lOsP0lHzP5ndmirLjohvIlQ
cwzsjrT2hxm+GyaFPrf3ZDBkK+BC2phjzPcgDnt9+PCb/OjBHnY4DSIoalFRXSt/
P0liuYQfTz4oPHeKNEWvygoAv9oVzVZv17oXKJou/9hsJVage1x2lY6k7F36aqjM
1GaqooZu5flJ+HkxVdQHcpuJN24HJLxuI067ua2dZHQ6A/zZjNsh2DxiiOzNn70T
2NM8k3zIQyxXfWnk8v9gh3ge/s56/UpsSk3dMaQ4exINwouQES8vCv0igCKumsMI
acftFqgJZxuLnps6TMvn994pf8hLb0sMHt2y7QjzTnrNpMPgqKNrp7Spr/tayriW
5DXlFnOu3ba0SEiUKuy/5WYFmdM7xdlb/8GKC+KwayTpDgChRrXkOliamW9EMc8N
nqwyhZI1d7S3PZySPg73dWsyEibfTvYCQ/LmOR1jSf9+Ok5jdGnWJlf4xscJ9iuU
5IuRaYoVXqaN81vn8Fmt+jSngyte4G8vOFtMUsyfobc3KI+fE2Wt7+GC5wSrbGu9
hdAScla40uET2wuBOPtNpqlSm7eqzjfLtEJKTLqdBorVl6Po1NDPJ/EWYgNxiy4l
n9uP/sAwbXgPftvS2vTNDj41NzD3aJtpuc84XrzkmUQWjVpu7T2AwnCiSHLd3sk7
bHGhjfsveznqS0Lq0k2EBVL9AV5FBd87uLm7GIfhkxKYJaSch14lAPovKeCrRyyU
BXXB5VaHIf8rGR/6K0noS+Sj6nvxcgUFMTGQB3DYwfI46qeZCoSh7Gax5WaNDA78
1d34ZRtBxbXVM3Ps5De1WtQtILGNCw0EthldNp2I+aR7DmFx9Zun5y8qdY2IYQ+Y
abgBK/r+H+VYIJ19eEp5mpAcSZ1SE2dKXXqJ4MoaQbKU8OHkWRPeiR3pHhRl2y0P
9uNmCG0q1m0vlWXoJD6FL26nDEEvzlBOPRYp758+3QhGjOJ6Hp6fMOHkWWFqNDov
Ud5wuGPdKO2+V5NszCxSz5fG9PUajtZKdJfMJkTz8Gy6IDu2jKk4JqCaBP+lx0Oi
QUbkGIASFVRjmyw2TL1NqA2cXwa41YuVfgQlyGmj0aY25H9K9GwKyENDQziL7SGH
kjvzj4GMQnsA+KBb3EFmcUST3tVkiqLXjT54n6S0r5k0uctw6Ha37cGLlyj0BPNA
qiC2rrHfDQyPAcXPUxh/A7gzvpjDo8y5qoMLtw0GTbB30Rf0WOYjspPdJmIRUjvF
ffA6qvYjdJRO2Uihp2c7JTg3Qr63rwScS3FLMJxEkaMrCjO5s3CaXKAPkbdEgq45
Cxu2d/dtVw10+2E7BJG0mwoPPxN3oDMnBi8ES5YDJR4vWjjD/2jBDPXTJGEWEiFJ
29YXWNTd0l0gtPyFb+qPBFecEI46PdcSb/zqSymn3/6YKbu54wZEexrQE5kBZJpF
FB7DHZw9/V/X7QCGdk0TEWMokjVNi9T35Nj/V2wVBYSZRaJx/YdPvtcy8LmQpbmn
WiAiPnt60s1Sryhhcp2GACPd75x4P3LbKf12/t/Ejttky+4G3SKN58hMktelfchP
HYG/827Ab3dCJ58MCoJZm0lnVRMtJiN1OfUc1NjOydGskW/W9YEw9zCof8a6zbW2
nOEU8L6PuXslc6c8TLYjAaqjR6vKoC6RzpPQs6ma9yHs5mcd+42CNXHrwUWLwD+G
E9T5vYkAKHmVoCoI1TiRwa9Yupd2BQwttAbSjbZtqPvBhPe2ooPa8EjVETr8vL5m
f7iW6V0l9hDVNeWDcYnJEZTDhCjOuwlJggB9hlcnX13SxZJB6NXkoQ8A4SZqF69k
Yq7L8jOhnr0onPselJqpPXAR4uzDVaTkHDU/FwG6iSpdFuV9Rd+kpwvcPLbxGhtI
ENjyaAmktCqArU06Qr2Hn+DvPs0TJqKwJEE3x9pwe7/+LYff8NjI/tfleofMpq+e
VvO4vV4koyP21gwdpBNPJNX3zJOXqTAliaqPcfKZoBX+TcXOZevE9IZIxQ/EcaXD
QrKme797orXa3NdYOb/g1bSYnDLg2D+RR5mZ499G9ECzh7Sgr385ZfCuSUkop7Xv
sPQ9xDgbX5Hy0PdTcOuQJMDIKDwSicpd5ocG8GzMf5gh4PPZb+bxLv17kSL1s+pR
EoRJ9QA8/dzrcZjBLbP1LL1P5pc7X6UC85mOFd7AVQwFuBeA5bIb1VYKP9i7Tpjp
+8K6xX6rx2vWdFyvx7b3pSQ+BZBX34HH81O0/i+9nob500raaiajE+jYJzcXeHpJ
Beyf1PjrbDrJYCgPduDA9y5+DCMkCNhxquPihsXjef9/4BriA8TCalhVr+EyDkPD
G9OPSLQba8bCLHk7C0nCa18pmtL3HiXQdxro7lmd8j/FRPkMuiUhaKleB6Na+EUt
qAfiRDAkH2Ci6WM4dHZzCer9GZguQhdF3gMpgAiO0s+oQsfajSa1sCXp6VyQ9k+1
5Rhg3sQlodr+cc3YEZ6LadcBozSSnma8qDfzjMreo6vTtPAWBEWugYC3pN2MRJBf
MlprkkXkhYrqULl+yzmo7tu0Ta9VwfTqpzcqlHvlduFBXFsP/wJVmpgn+JFcacgF
RqjfDK6jpr8U5YAIX5fIbYWTFY0Ff4e2cVbhf3Fl3V/8aLCqTC1qJ8X1d88bmyV2
m4iCs7UA2cGQVrO1ol7Xlhh79lXbNNOvi+FNsJnjWIWtmc3ssacdLU/wMQ8ljRCO
BVlN+uUz3eoirQCJYr3eAyHF7QXqZ6ziU563E0UxpkPxvrn/ZzVH30resY1FiJow
i2TY9if3HhWMknEKRDfJk6kta6u4Fw12P702zii49MI1kzs1qXywuPTUf4dqh+Vh
Gn8shVahnWyKzhVRA45sTsvul2rLPn7OzpjQsj+W1uftyiw9BgIjsKWWxdoa5Ub9
UA4b+7FCO8+jV66u6DbWX3fLj5upsKXhO5bVaxQnv4rQJsiCbKSe0jHbUYSQDCPe
e/zLhtlAqnrF/DacxHYSuLN5yXu6+yyZDstzdzwyZkGBAQHF5QcOZhm4M/K4SofC
Q5yJoFQb/0rFcikzoIV2/jEBtscf2j0PJ2Db4iAujyrv4FvV/lcRyUNSIBCHLMm+
gDUj+QBozvAy3CMksQt/jo03pwhC44eAy090wwlFhnqDpZaYxaslnzEJyngS/fUO
XTt67oFZyOkwQ6p8vnMZ/KI09FK7f9IcJ/E2vEmgXcqIX8OsdncbMVKngak1mn5w
Sfk0rEkYy6VTye0T9WbSBC7XowsEL/cSz8qLNTP9WVlOdJObbYXF1Fmd920EkoHL
KYdWmoGyaCIfhRHtlPw2ZO5bBmlCYYDAiHRwfqJaQnpzbVbDk8x1cO5PQnS+4PGC
6bnCjFofwrz8yMrK10G89PfLyuAb9CZVG4gj+EhYNJCXLiAjwYFav6MnGi7mK6H2
l8tLhenCehAyt8jvvTRpRAtbA3cWHJI3IdkhnlqLKt6u7hZs2Pga1aOVzpd6SJSy
F0cWFsrdcJ5B0RxwsYz9rJ1hsqqTifiibfuOJWEXopJKd7CevqAXW3sx/bdYGLff
Pu7ZYjXg1JBrcirML/DQa30nQQAY/qrD3nSwFDfkfsDiDxxPHJ4TFIxwnD3Hdojv
AOvd/t298KT3lD4fhX7FKjFqW5k714rL+ZfRQdNwEQSLF8tDQpE21kDC1TquA1hm
YA/dOWRUF8JwS9K21MyPAMbxX0YZvQ3xWhFC9DulyP6y3gTPMjyyEccXt14I/zlU
fqE0q/TB6L6u6WhHAZoQhvb+Kh4GiKcg+DR625e26/QiK6Pz2JDUOvSqZDx9u4j8
3am7d5No4GLry4AarCLAzkjuVoT3ZpK37Atdbo96A0i0ckWOY/w5smWmxbSgn4bm
RQxcF616PuYo0dRTHalcmJiXfHRJiaR89YGSjUb6I99yUf2oOIv2xCaCJTtvzB3+
VT4C+3r8kND8TD2ODn0Oot5NikiV/4NLJdAXKgGqbiB3kErHWgJ7mvEMLaiPxJsg
BwyIlNttryvDIDYIc4CHryErl8EF6wil05h+6kph8+G+98ArCORoTVRXcTJ8GXfb
00jkwi9mNN3OZ2KXNixEbHb+9WfamZa5K6YidODVM07WK9HrK2nwcguA3dMhWpVz
dqzOv/XyJNn3G8hli0xMsyneX7NR64VEER7guQptXMsH79QwsZmZfohcJVrBJ8qJ
fQ3BTs5DKEGaZ8DFt1XevhKSYuaD+YiIgihJc/yny7zr6pSlaXV4ELcOEl9z//qI
t/hlyPMlt1Xi70ZGi3nHaB8LcDSqmkUv8cXO/Mb9ePbwxHoNBBUvsqywil+nrRdA
NUrBwgT3QIh00/HPoL3UZ437aHEWq1L9JkN8vTR7oIZwim8noROhUFNkLLHOU+A3
hr19mtjsdMYML7q7oNdgcvsY9gk1TUzNr4/HDLy9xUkLDoTArUubi/D+yA0l9dLq
btsUdoX0KsEeh+vr2fvijmDRrIpBkGWbvVpknNS6uGIGvk3EPttVdtAKd0hUMgco
fDpwaSaiDj1eDtL3KexzqnK+XU7mM1bmERs4lPoIg8IvPvgy09qp472u8/48G3XS
bFakwdkfDqouoeq1NyIPcVzKNRdHVxBypXlT+MVrOwjn8aVjivKn3e/bfWCERmlJ
Xd/S1zTs6g18VKt9EpIElGvGWUiEg54J+5W4xfrdf/Nw5J02P6mr7QkvNm9iUo5F
5s/pye0tkThIGLz6LPK99Dktk3C6+qW1INI58Od3sUjXzmotwboYibgzGAjtrYkv
Gj9MXUn3m/A0SvtkTPJCQLZkhJAeBgy6klZMJVhzO9BXdiflPPECP5BHAhlcjIQq
pqFjPraOhfdKPEF7LYEDlfCejR/NPeWrjZX0szVz2lM8J8/XrrfvEXzIhKGLMgRL
NLz9VIxRYcPE7zhiW+f/SzEw8b/qPiOtDyW1gMjd/CYqrNzFFQwv3UpuBBy6v7lD
iJ47w8mt+KgV1366fyVpfnpXpuvIseDvAZiXoUVVGipKMwNcUMmZlA3gsBr6Io2k
G+43n7cq0+97MQx7GtiedLBuFAUJJWa52iTZE4M3xs2mU6xf7BafvgEvyYiErbn7
X9kadcBJFMZ3yFLIEyVE8yzitwZ4ceo57OcxqFCnJeIyhWsrw0LgqgMVL4IE5AcN
doUrc7ynsVTkDt/UOfM4dmobZOOVhcHfPFEZysd7gwkV4fTk6H4PA6fGPHh63dO4
LxcA+gbqJk6b94QwKUaCmtxi864nLV1DegkxNxlA4iyCiED4VA/g/i+SsF55CrTP
ThNcf89jX1UMNc+FMX7jMSH91Bj6ILP5gUQ4nHluU/YmFX76Qu2haCR93mA8mJ/E
119jdga/SAwpXdOw0J16hEyAdljs+xh88BsPOPn2tAT6ReSIy4JhlX3Soym2Ookw
E6iclKmry+oiuIbJJNmBfeoxaNQ7345Wt3eG76RCdLovFlyPWQHPvpC+PDgTq2MQ
+BBfemMaLrUAcHC9pQOy/uORPzAqPDHGQG0FAqKU8n+NnMuLSXkS/SPBJvM+06Tk
toOYqp6XUdZd+cWNAUllVvMiCpB4jviQgoW13z/dzjiZ5hjZYasrTjIJaZklKtAG
l9J4qH9N/MszPg+O7kZ2d2zDptTLkTmrtOWnugwSfVr0zfsf5jKwbwR+yo5kxQ5d
5N15wX3N/x2ekVOwlNiraOnBde6K/h0ToCUP8sXQmAgVbcYP9Fl+Ji952zf0k82k
etSF4jeiIgLWJc5iOBtesnYaoCi6fDwjMx1bROd/OmVCHD9y3QnMjTrlDoSRYvaZ
xzSbgkI+RTp/tAEj54GRtsQYNGSwDQ6LWZhQu40S6ssFUNt4d+hObEHttn6RBsGx
21bbOaRYeES+tqvEW1McDvSoPSdkXcUn51MaZ3x+UqHKnaTU5hFJKUoPYty1mdD5
dkZ4iXk6LKh6KCMucRsclDUXNRjpB0uIsA7wL6viAdC8vLwT0ZzhIKniPrCtS/mQ
nwl3+hopuhmNzMVC4vZOjoMTraR8vX71fnEHrVL/50RsxcIP3neFJlvYNkv6YTFz
wJs93m1kkXRgmr/HRrXEoakG88/QCySTwS+U+uk4l3EifaVBOEG1Oe+jUIPjsZI/
ulB5exvNuthX8yAlX02Y1mBafWeLVNis3PbZKgDHinYwx5+WtQTxgSl4Ethq8fJK
dPpF57bq22YzaGqkWofHMWHa0HpZOePv/1GntJC33dPwvhEOHfL7BNEAaARf+t/v
HpuK6TrpySYav/bPu4kEg2YMXTrqpG45lBJkVDt9RTmjFb+KMpSqi4Zpx7acF/DU
tFJ7i2z98hiSbeNksTgS8wkGTOfrttL1IEietPgUpxBScoMPraL9oi2kR8Py8Ul7
fU+FS7T2N0ky2YeY00lcHv244Tdflv+Kqsbze23bLEpxiD9rCyd6gmnGOTlwmAzT
hqeNDrGd6ddOReRv/JnXVqsx9rFzNvprtbV1VOr+/5UAdCdYSaUKvSe8dx9dXcSf
wM6u5Ffvh5ddqxs1rXYrsngLqRV/xlgH0jWtYGGis6LgzfosKVcoVwyjd1I4856t
C8KAgSLLiUjMnIowhBensYQ1/KGtQ93w8sn5scTWTogRyGMJh77MJcbGwGxCTaWq
G8kgcDUcH1DNSZr73+HcDfRxnJ6Hs2jYHnYw/LOiuIqafW0zx+gfdadxKzkcNqmA
6NHPqF9yJkajNewjVkIN0CdIt1xXh/sbBoqOez5lzNtA7UI2jSqG3V5nIhvtGbp1
ihqFPXadtStMZLyUgUGz735Ie5toPItKtCZYPBiYuXgMTBpTLOLiaA6PYNjbUH8N
EKnhQJXujiXI7oD8658lrdNVaSB6IMHopyppbt7tPoux/A4Dq8KLAfH/28RmXEwR
79ErTD8w3HlIbruXtLDsKR+iVKHqbmhReWZBnGj+8eI7AUKtzvsJL71lzs3k1SOt
yiOmFWPjKougk0ydE8XM8/Zha09oFXaL59qqzL/rUaOpO6/0dn6+oWHSmNpz27PV
0y/FzqR4GWCpiLvHTvZdjDlJgby3ymqHx2MvuB36SI3inqrlRd0gikCQwe8Ju3k3
eIsVHr5EjK7O4eq4f9Jbfh7j/DhJOkMShoVRgAlEAEL7XQwJOfOPETTNTh33w2sl
LE5eG25gB/glgGTJ1HjiiS/u35m/j2Agcpd8Yc6b7U6jbEdaAwsZMLLr/yfGZIZx
qpRuP7L4zB4COlyP1m5A6dLegu9lknOeFeC5jgp33l70hypeAcvu7lUVCHeUxcKv
GZ+WkK8yhkI8CGI73ksB5grFJtg2gXrxLbnDXMwP+If7mfQX7ARFCcCepJ6s2Vvh
T4vCfcCjnr2hW8/+XyMi5skAiFM8/pJ8nL0RNcQZlIeksarNpnuSbPH3OQzEvs4h
WZxhW/de2Kzsb7jv7Z/xLITTytcMLZWEz5Vhld526lSVERYbR9u6uOCzD47XIXqg
3xwn3p484cmZI2lRKS0zk0LNd3IIml7MlJN1xOheKtQYGiRw0tEkYzCmBv4n3mo+
e1WREtV4zwIGQR0iobz/PfwLKrRO3fKrXOhg+43h4JxKQtXIevyNiB+5dDGzeQRO
vecfZkUr89ciY0dpfX3ySs1fLDlmIrdjY6KbtewcXlh/IWO3t7LeqaNouwK4tVAj
enAqwJq/2g+BPHxUnw6PzkChHnH6OA3IT1drnWg03e2EmrrJVJ+eSdkbkGn0gCtP
uYA6YmkF7lLyY5aJcpgtTpFyEKP60R7izVdSaT3R7mJOeUI65qHB9VtEGVrkPWBg
dHU/nhhuQa+wkJC5LZLbdeiewZfZdWDucgqdAHU5f1YSJzhZdRC3s4bczPT77OdF
IGJ1GlHIRfEVGNDCqePFx/lc3ASiAnJID0kjkepXG8vahkOROMaLI+MTzWBBu0l1
ixZZY5Pu/OEoO1lpoVW8sILi+thK6FCCYwa1svnOz5jeFOXn/nxXfHc6gx77xnfu
ElFdHOLA8N15FVBLSyrJ/jVZqaZCfAT4SSY4UUE+GHheaQJNG247O0BX4dEoc6yC
ZTseFEKfbHopCXdGi3UoHgV/FWcirKSlrfFtKuk4JHObuA4/n+wSAfd7S6sG7GVz
bl9w7RosJrt9SCAZ8Rt3M9ccq0dz08apJgAAaZ0w6jSrYDL6Sy02EtXwBjNvROcm
bu5/aV3qy6l9TMbYFtExzR+Skkd16m04hu9Dz2z7L2mE5RH936oxQWu7+LKEigCO
oeemIlOT6Zdny1v07Us5b23IuSVfKHa+j1oEl3+0FmGPxlbFWCP8ZE/9YiO7M6BF
B8OdzpRKBrr6CWdCbSHrwRh4HxfLj+3EVF+RxhYdzwTFTfCcsjKUweRmB6hcDFqd
qAMu+YAfN84C3opX7cnhI3rqhUkekhgkl+WiKEnZ4ODgALizea1AOi1SAH/LiN0+
sh0qolOY9P/hbZzta3uLTw59LzPW/vA6azvh25Tx93GJk3QZtM4EEi0qShAGZ5dC
j6DvVlscYEWfgvDfeUCctl08Th4WZuW4ZJn5Hkv0xZ5oRJfcRdInaKQg+QL14k32
RGqw2Ubq+7nsk75tnPbUCSjffweWVvnOzYyIWDu/iTWmLNt328b+gthbhfLizvGw
LA2J23HNjyNHoWaPJHKiDyNOeW16KM4ZATASD/MINFBD84hM2FpOfvIGz40US/WW
Xv+uEO0RBl/rHT95A8Mn5bBrQrCcXtPO2C7ztBxBWKvAWMxPCAChVxn//fVeoHnc
Y/m6u5QIB8bUBdvKBvYEhaONAqLzFfZ/TwFilFnUjJfHjKOMkOsNoW32TvfPboa0
dp76tPgZdk8ucbyE8cqh1F1ve6ZZKnXX5wKiFMeewv0QUDrFMvhQt1I9h9i3ZNdj
4NNkFD5mgcfkd4OHMzaS6gdk5MDAMbwGj6Cln2IRC/47uid+cNrT90zzr0VLSNSK
EsXkva0Kw5tV0/J5U/EGjJiwFTqgPbcIs0Kzp9RvARmB/iFhGrPsuDRMd37Qq+xQ
1k6IRy/DpXldigbTy1Md3EqWlIjio5GWRfTIV8hW+EPSkCDk08paBYObihENmeU6
EYGYxDu8jZvCaRw+ifgh8z02wa54T/zs8Pm1nM4eA77X6ayxcoVDEcvszOCcAFaq
1e/h8XOZiGY1o1HF070d2K7Ktl2fpAfdVkAz0s389706+ksI5Zf/7NVFr5CEcYbO
8cweiVXq1KWQopQzXNTz7P0ee47eicpcoF7UKQpsdhV99zo18lVwb1JwV7AMpYWz
hX+N3b5AcGwe5q3LAAYpPSK6Emo0wMS0NcDlfk6OWp8+JaNLSU9fm7GZcuk+d5nA
iFmTm99d6tTF+pQLYVZKGEgJ2yQ1MfbiWwT7gChBeobBWlNr2Q/k1BniAsUOmXI7
PVG+LDBIV0rk4VfBv4SELADiq1f6Afslb5iGLhHoNTQTv++l6ZoWqKueaUn6yc1k
TJxbEH5cN+v3HYrfjl1cH3vBrWZuCdiVRGQf+F5C+yTZQlE2yb2BqaKikm+1t7iZ
7FdHYrEycViFZ530hNPar/mi0LvlRMRFujQwQB2Mds8JzBpMaXcslq3Cc9OvyZgR
otZ5PLZUgGunUYsRCGl/JxMF8yVcXKjZxhEN794z4EDtxFi3nvhmJb6JdGiPoi4N
2TMX/LTxgVi9z56Eia+P1zAsZW8ncKdv44EXuB2RRhywtPJMvZeuMABez8I1+hhn
5tP1p7yKLu5Bi/qBJ4Tu6RhjxeLa7zlsq8nMv27+GsWd/BjDhrrB51zylkBL4ZrH
buKsTAJzzB1Dly1Rd7YzjQdkDS7Tqex/ZwdUnE2T2XgTG3gxOo7mB2AG+wMqTXQU
oEpxukb8FCRlgG1+kvShl8OZvLAzRLFIWx8t9ssayJRs+4VxKdeKBqI4BIYjW7GD
KkkyJVnqGPTzKZjyB+8mBx5LvsSrrJ5wULRHyFJnY9ryg0EEVn2jsjjd+PrOtMj/
ZddQdNzAxU2sRk+u/+5QEGbJdQpkt+fewxPSoBkGOd531XSR+bVArtE83c3g/BDr
EwrZJQcKOwyQCyA2iqQCZckAyMdY0kaOU/xUR5ZUpqz/ypD01LW17I3Sc61ne7Vi
Z/bQzTc4jA/+Ese4CxuBr2y2NDmwOkqflm9TogNqn0VLh0iOAuCs+96AxyklWL4P
6ixGeCx3A+vtpD0HEzbmx/E2klB15utdl59PkU2tCAbzV/wgoHjMQFlLfbg0guno
7kfyJ51VZGER/R2EIzWHMDYaKe0XFecGl7XoERIcEDy7PsWXpiPUC1MmX7LQ6Q3y
k5Xy8QCw9GoT6Le4UOARthzW6G/Qz2hppbvfnZRQvn9y6ZyZ/LRoL86uP5kK+ByJ
OC/oMW81kW65YtqYl6p1RcgyB9kj2Gu8+3CJDDtEytlvCC9zygRRP7HyeYGJTf/k
3mp/ohXSH7dwGSTry5Jen/JOgYAMCpIuMbVRU5klJUMQGXwjdU4+jSBGCAuGRcWJ
uhLC5xgjwqZcxPXWOkV6/PUGgwyisl0NIuTzGSpr5KYBdLiEtDOf9pZl+ZMVBq9W
LLPhJmkCvUJhAJmSiA9cZzKgLjF2dS/VUvFMtYwAGv5nXOZ1Ba+tBjMvHm/EHXoV
/A4BUWjHOy2Bs3Z3eG+tlcDZ00RJKnFGvRQeXeEv5MDeJw/ALwDrJd9qvVWdm9TO
5ULq0u16+NvspGFqGcojozt3F6GXqlYtZgTbnWvzoxPnB9niYfPl2jftleqO5UU6
hhVmuoc4PpRauLVY1XfpqsREiY6MHk5wvbvdd+LL8zAWYgMOH7YnxsaeJfIXfV9N
0+8D7C0aq20aECCpLu5EdkDcAP4Z3+ATh+A6F36clS18aEHJOXmdABYIKaM5TCfQ
o8gBIV8zy7rCFSlqbLXweYiLuTEmLvyR0g9318dJyulq/UDc/JY9bUdlO89kIo7w
bPk6Z6W+UQv5XhbAtsXxO1xAHf4whle+PNDgiVQUoUu8iG0OvAvUtdw5ZTwukQZO
i3MhTcr7qEYpZzIvigjKy6Z2WpquTjyyX3ySxxf1mgonw++ESBVttfpZks/RL57W
qhUKsKl56UVB2ZvUzaY42edQluCk22lFSR8KjB6+T0GVcAsSamCogcwUySKaZ+sv
5myNCEz56BKgtCykx3D8yiJEJ5bFmT6aWJdqEskGqnjmRus1ydD2RSIWC7rTqkg0
AaldlMW9r2Ff23vIs5QvFB87W6fjN6UkYUPLRH4wvIkd/keRmSPweP7sCLMk/hn5
x0EzW4ofQfYLCA6umfbRD6Z4nTQvlXcrb+S7yiM08lB0bOhExUEtZsYbAARJ+K8j
RnCxUkiTyIgon7yu69ScnbnooxSXf/bPBa99D4AuJDe1QDvG8/Nj96C8/X2M+hxZ
ly6SC3UoSrLxT4fFPc0coiiFz3YdD9p6KlHEQutkQURDjX02vLFgXXxnO4JJwQLh
OUvI+pY4SkEiTvT5TfIfWzq586RO3GVrf5LATGwwaA7qephLmJmdJzTMB4tvOx6m
5AxDgc+Wjd2rrDwRObsmp57gubfQH0Ih4Dtos4JqS5Ai77klIVaeFet2F2yON1iL
HLQrP35qK9/eZllZ0x4Fv/Gu+6SmWN+2B07ke/4ABIN/3EHmUAAPnrbAo8jrbnN0
eBr4yyNO6z2beq9PgE/rHKIFlavi1j4EDb4MTzcHZQWeEN4cXb+L3+PC5drorg3p
Gag5a8zKRCwDruO3ds9gep+PRYOucfZri5Np92WkTpB41S5PogEiUpDHt01TtlUB
CQewSSn1zA1T+8VwJD7wvWOE3mr8px3WSgIan4tNAZKWN1FUiNpCLwFGKkr+ZZLb
L7mdUI8RPZSLiUhy/ZPciGIfXomuMFIIayV0iQndJAxCxnod5BXSMqSJ+kL2xc8l
a8kfrh6vC9nFSgTmx6n7l+Lj7InU7MrcFNKgNgCWC7tFE58tpVyK8sZ6yxlL+hm3
4Idhnyn7DMyjkwB+sgXwh9vEsme61EuV0amVU9hTwlOiaW267Zn294PJWqZeVsw1
ehu0Yzx3CPbC4jeFoopMjZjYe8BOZj7KSEPX1ZrX2E7XZpJ02aA7AX7IyxT5MElM
jkNUJ7k6iU9cqmdQcSbIyIthNymVDORUiUP67k/P+rnqn7VQk/kIBq1y57bNp/3V
lIOZcACFzlrGv8Xg7Qi3tLjt4jCCmMtbn6JbdIylXjHwDjiGnTloCNl7Z6HCWwNx
9Y/+AK2FTpsXScuk2XGLeLISDqcAikwWAcd2MB/7sxIZtmBON51EQ8fgLrJGrDl9
QDtB6M0MwIHsSdJwNwV/5L3Y+FS8PQMCwZg6egB5l/+5qFELgXLU9pCEV2LneLDr
1yqhow8Y/Jsr9ejwABjrdSgkroRZjZack8S6v8WYQegJBr6qsG7CvhnybvCM3Ax9
5Vvzua54+fWnoaCFebHANqoiNSxD+9vX91nr69eGa4TX6a4zqcg4ZlVj5SvMiuFa
0XMmymp0YiLU5vkS7EEzde85iUq25A4kZItvCkJeiAmvZ+UzmFkEQNfG5eE5XfzV
TZcW0tvTXUo3JFuuT9BMvduzWLAE9ii9Wyw+Z4Bb7Y5u1LwtlQjNFy1Kw7QUEDqm
D51PwYMkmJnmT4tncuIxw64NQTSV5aUwNNWEWw/y28AT5uIDnkN/UZEbThpZaJrX
A1QP3lS6FszDU8CZfKx0oy7hlq5Fmf7TGfpaokaI0DRo8Xwxah6OjlotcyBdnnIM
oljfSt4wJr0leKy+AKgJBFYg7REYm+IEOfO54hVXjkUO4IrQiF9vTZ7jLzostxHX
KcBLeiiVmgAEzXlMKW7LsEGbMYnu7FWkyoCt727Dv1AOeQoxv3LLBeDdLMSVYvXR
2BwsYMnpK7Qbsx8rQKzpS8ewiy9lNCGBZxURviTuNjar0pM0GPV8xxBnyZ74CtRS
n9p8DTQvWnLbn5lfVRqM51It3aQCURLnDLTeG3DhiM4Ye/2itFXMfGW+tz4obaVr
UgjaWNJR1P6nZGubNflXvEU4a/fx19rKP1Jl73ATmvyPcTjeg87cm5VLg4/bEeKS
g6fYXNkkewuTzHjITcFfNxZmONjp/HR5uSqBgj9DK0HrhsqmDNL7Boi6r+H4IPe2
k1mhVa6yem275WHP38Z8gRB2XY33ZSk3WTLDtbKKRYidZKa2mFsesHn85N02aMiJ
pSsE38vDCN+Rd74EHeSSbdSsdZFamgNeUQq71jvlwBoKeJnPVLdTP4aRnsYyhPwT
byXqN656/q3iQnM2QvEEc4pNflLtXI9F1IrYOmtdIMOcd0MYLOz+KyouVWwLwg3z
bcsF2yZCQLU18N5u0hwxONW8z2+dnGi8z4/TCliL1l90P7HPYhcgEZAKEnxNEiqJ
Hl8BwkOGPfRsT6K3qtFCAEO1AV6XwDHjOPYmCbVvvx6bSXy1bKNsUvoBoqiin4V1
dfWs9hkgHtbOq1Um5fZIaq8jizpmKSfT3hMfuzqugfgvr8XykFIiLdiJCOUmp5yE
YmTHCJfOfCot/Xn16Ut7EeDmCZprwp1SzrHkmhZVROkmM2Vah/cX18tyd3SqhXtP
5wC7AqatFYjstAypDSz4zO7yj1BxpJPmRhGnJP09x+8TDPZOiMIcnwv+0PeWEt3o
6mrTVCQRpXZ0VWqNrbZB/2YE7A6Ubq3uKrS9pyC59xS2NCIh0HqT8AYayV/bm8m7
/USZSLyhZuhSy3KPRl3UkVnCDTIlPjh2uSFqq0ddXhasceJkBmv2v8nuOzdk0x/w
3Ipl5+b0vBoaLOrFZSFIlsPg7YtIFfkm7rLS0klTv8yRnALwvat2af7pA8vmmsbi
6XoWSLGhZQPVMlhL2nfvcwyF9oIPYU5jevqmztx1Cc9sApHrlR6kJef5r2eFIeJZ
hlovwAjze1ZB2PCPCngmG1NNMBhu3yDY6bRUKj6610q79bJGpVTkYiILUC6cDcvw
HwvnuDlA7CyG5VEqYZsNLlaVOrjVWprVhge43UTFkyRXiOyp1ZXCg5lkyDA4Mte6
ffhyVeqy6R7FBxbl4akua1nQxxDsmnmtBWnRKmXkIeM5l8y2aPXTRqzlbsy7MdVu
Cby5Thh73USFJ/OAN+lSeZoGT5X0/fq9gkdQW81SvfmT+b4/Sjvj4O5Wo0zLuLOR
3wZOUMlunElL4JH8ejwL6W/bVSzjunpBG3k0VbeLNbM1c2ISVTzlZweHvwuivhUW
Y5NSFxh9ZBcDyvBpmjbqsFMB5Eb0Aj6Bl5GR/NEl0mQ46EcF58vxChv43kKlGmF7
h63+zVhLq6vTo0AD74uS6GMwjp+5IW6Dl7h/EY17qJzg7NFSNyPx4iVj2NUKPvS4
dMgqyNkt6CeoWg0GLE2N6ahwYFfuQCPhKU5rp7OCi/Veugy1xcG134bydmgGcNvg
U9U7rEbtxNivWiOsa/bUVgzDXYveBcZV8K+ZocTKzZ+CXzCPZjuc8NLa2bHn/XbY
QSvTAZOMzz6vI18LnLAZcL8BprrgIF67dUvEnSfvov49clurq1vSZiVCy6zjEg6g
FZXPl/OxA7t71KKGZQOp2SYdRStbs4bvxxEFM2O9QbGMeCEBA6bKQ5ffHcdSqVew
DDZwuYEC/1JfDyNk3bbUfW3wMrHOk3j7//ekatKt6x9MUeNJs5Nr0QW9DcLQ31p0
49eTP/YTcxbZkE5Rn8pbgJwE3ERgfYcM+PdDSacAEOWdx80dRrIZoVMC+loWppCT
lVDfxSN5w+71XPcVkhCKPdlyl2B6jP19bKKgy8YTmY0R8qOYhvuF1afsa0APrhZ4
oV0N3EvcBmajdzCrSwBmyeWWPH2SFV49JbETKVPa1W6dhxP+6HsA7F5LQ/w9LmXi
x5bNJe9DU1B2w8SYrUIr0asnAjeYJC8DObcKg4Nb0csGCBrHJzzS7iIss2LfNWq4
yX19fAihb+ZKdjuLIullhI+Jmc1+l3tU4Ls6PyfvGrTXAjS1xiMNfVsCmQAMYhk/
cn51th9SOf45CxYACTt7GguocBi0NVUYYe5q/U17XjCByTWC/ME1p7VEwy+QsNmT
fl5VT1FvH6Swmj4DEe/tpRh3QZEAEELLupClyDP4ExPLhKjj9zAEwRYyKuPc6Okr
qcH5qh/eIodAJODtBXvwvknMrdN13PyUnpeO9eS0be28n7KwLXlPwyEhjeEi0rWY
GGpDIVDe+Y8YMgdEQLOmoJRcvdzwTd22nOPGI2RkqnOSI1c5eSD4v+60uapsW2+7
9+JvDRF26rBsXylk98m94zUPr0O4Mk3utbFKrBR2PwqHgsQe0VI19rEnIJKm8Si7
gZ6tnO3GMZ/yVkDSXlUWDCPwnMR/JxohQN3/tSd5LYaKS0LVoyahj+NUOebts2BF
Mko+0+9Z00FpJ688a74RD+2sVRaHHl2lVknH1MyLb+i3FJ07c3f9IvlIODi1yoJj
o6vn4Hs5O0JZdc7B/GcVNOtI+4TU8FzgdItO3lnSUcRvmEnHWFHFwFl6ZaozPnPQ
RdVIyymdxh3Q2HQ5/7kCNVdnQueYdnW9hx3cIDSS2EwbP7c9T11BuN+pWajGd7Mc
obI3Y+cy5iIb3xKfli/HSJMkrlqsqA7wxLq583gmlkzsXgHCo+hnxIh4UxO17jYg
s8Pu77HZzIzaCb1sQH+0ahCCiSKXwxzu0X46mt7ys4k9fV1N8SNFHpMJnpyj8UTI
VL66zDokX0y7pzuLHnE/gSdBBfRcmODmmum4YoJJQ5TEV2gn0a1xXNlZKi4ah3F4
Zz/HkRPZTRRJAlhjsr4nlWRdQlAcEb1LyKZenvhFloe61AhLwiQCMU5H6JDxovlH
7qihJ60TznmsIf0jreJIJaHnAy44ufAcx6o/jn7+EMqT9/v8lsQJQosJVFbnfspo
uN/aokZ0NNlaB2lzIGPBT9orwbHDYXOFXfH37PWOjMviYmMOXmqlkbuM5ivXaMSa
d+mQh5CMrdegkHpwC7510DKCH+ARf67GEwqG6WXzoCyWtIDi84JVFlJWAqKyoWvz
5qxiucMsLxcKqdngLaYa28yTy894rMR7jmJTAz92XiZukBfcDhHPwaPELXAaGIEw
ir8X25VSgNWKX4lUxX7wSVI3z5VDP5ls9vPCoDSh1o0gxqTDZWqtBq68EXOptZyy
S3EIfh49rbcE+3H6iPiQDw/Hk442Q/5cxTL7VGoVRo82JzLteIT+d6LAwit7T8F1
ozqa3CWNsMThaTB4bL/SWu+xxxP3oxsoAZ7iwIztvbfM14uM+laHXT8xeOD3lUQB
7bVUFrzl6TVvrn861dx5ORFdG3rA3nXu76wh83dEskns5MC8Yul0UPsYpaGgGedX
Xkg330sI2YGkdhBv25Xwc5GqTo/Bbsl6VmnYIwfszlFbQJ6QUvtxhsrTOTc64Kym
efI8SkH/Rm841GFf7sgSuzjx2fX6QJwKDTWs+cwHME9udqTGNDF2MwqU9J9HjnzX
HyVSYc9LBVJOT2U28C1K6hQz2jRP7mUfzMUlzaYB6OwOQfMtNqydqGhCRIHb73pg
RT5/oPJD28jNx9H9GYw/tU7r9Rd4Xx7wKVs7+E/5aQFL9zOHHBTSzodA7YvXIcIG
es0FUeqO7hCVJ43j8gP2wJOB7eNr/jF8Ybz2pvURpfjeoWWYLGhtpyXm/ufgZx1b
EwGmIJBBH/h2zox9Fph3arILOFrD0tSUEpfNqcvFM/KyaXIz+2F4wZUAMXsoF64f
IQ4MtOA6E3tJpC3mU78y45U/gpo39wdrlAWoTJe3JoP8U0R/OS3bWfyov2PVCq15
D64V3gUoqcKJ2i02/5EOFMSSW4eXcIEea6rQbHf/Vmpz5PmgPJSapJO/O8+jefQ0
Kcu8ITBpiXVESB3aPXlOMpdQnPRA+LSFF3W29kRZlHZIjBYzZwismM5EdQo5587t
IepHGYP627NcogDjfT/yR8pE741MFh4q4tp96biS6RlzlLjZ5tlmgBjje8nyUF1p
/oVaglkydTE8koZGwxFuTP6oon53FbLTSWZ38vuQ9UOFaUOKJ0XG2xkWSCa/bBTJ
+0wMI3LV5NL5k2I3jAS0rqw0/afDW+phIrOgW5HR9TU1/DSeUT/dO5ek6GL0nRG3
tCH9/9cp+3NAQPuj4yZM7WN9sBbnO9i48V3Jd7htMO5r+dbULts2+L06wTUQnYxm
WF2i5FDK5cfFgWW0Yhjf9oQbijzz8me9Vjrgo/h9DHKA272EzHDt02lKkXZkaINQ
o2kWocgFKXrbJA56OZiKBRKQ5ZXri+lnjt4yJgKGJ2x7weGeIQrN3TpHmb1oQqA2
TUKuBFSPjkdwGthG2ElYOzGmPrcCZJHMcA1kz2rVSuAYnLvXxqSyuHVkWvrrt/aR
HfCQ0ghRWnRA3eHaz6O0cGIgueZoGABlON+WC/23wc0W0NIJnn2JbrU9GBivfRlB
zO+NpSoFJ2Je7WVlcF4z6jLGK7e0Fkf+Ur/sKKHiWFPVFMhwjZCj47Wy4wzi4BIr
4ybNB/oTCG+0mtNFL3vsNq+Y4hqeul8DwF+EDaTwnpo26cZLyncSR7SmVK0gs8UE
rTxwGP47ld6M2HOfnn1Hcne10EJ1G8BraKv/nUnS2P5glCKBCKPWCZcdF+bbhV/Y
U0+LB3sOQvtpUwYpxlUuqR15LuguM80VUV+bJXypVvNFkfLW6s5NE1oQW0CuuK0X
wcJpPFMC9qIkfF6FQPmbvdYCpPSDG+mvEtwX99k1peN7fC/hjyBF3BfWcJJpRr+D
IJekX0TERKeG0NC6k3+mRbrqaobujuLbNK9xsuXhFbHKK4ETFGILqx93FHMcilRK
qXL4VPEkWlyB6QUHrRUAL3McTil9F14YK4CORFQslMlHe1FqKNTTcftXryjfCv2N
OwA64kitJUmup+ifoMiysN/qKiPmGfJ+JzNMgKDGAmX4IZkJLyzc3n63sG1938tj
L73ADn5T3Y8iV6C3C0IkSglppadPjWwO9fKyLkpwCFEZf9ixjqeOgfZ6jJtXFlz2
+TPdnXtQzvlU/CmpVfaU65MpwAv8SIai58GOrbHagnn7bMVoZOMQWEeBHugHo1Ub
lxstNNLfUt8VAW06QxdLh1uB3L0gRjuhTx7286kkv32AQ4ri11ch765DFX3mk2wu
ymP7iZUHsmOe9LZ3ZsNS3CSoP4p4oOxU0F6j18YrnANyBuO0/UQKOVub9vqJOqbz
B1MV9e7NjXeVX/uykdbrXpOzxUBrNXQv23molkdDRsNA2pWGyO18ShXtlqaP53w0
LUf+GlbQfZVcHOfjiQzPKNz/X8se/jyXmVtHd48bbgcw3Qpkg3SAL0/ZnPQsAxdD
ArhkEbXDZGIky/Ya6wd80z+9gqNKCMZsLN5auyn13Ey1E/B7eIiBiESY4NHP5/5b
6OS0malMBPCGcGSPGgS1y6rYvdYkGEnhbOewBzDAnLT/74tvPI1JCQU+ozKWUeBx
Lpz0LMH9J62ZSWBt+/j0CKXFGfAFc40ZSR0Ha1XgIy9rjmP/8t7QXKU6hFeV50xF
Ny64ttW4bqpHnMX0tWl+pL4wTSGqRTTbMeoDQmhh4S1IvFnJMLOLyoZzpViYn+27
YuvK4K/N9/9p9a6DKtv9mM9jA0kBsD+AJYqTqw9F6Gnb6beWM5yzAA4ibULpbOf1
bXWZfCafFzTGRMdqwtwb8Tn7TvEO8W5uO85fBqZiknv9K/Y2cr/sf7YTzcYNq4YY
q43HZavH/TSDkV3JW6nluaVvrSBwOciOw+oCPjOMNrFbBFiO9g/vRhJLpi9peFQ2
Gqlwsa/3/Kgb2+nV0VBOfDh1miB7Vv0O3ZecZJ+P16ePFUfvoLV5yKfU4sxXytUM
pgablZx7mfCv4BVfP2bJbNZOmoeQ1U02VgVt2FJhX5k456CAR+gwRwSeFVG/IOjA
54b8lNkKCXTU7cbTrVcBUb27PaDgIqPZZtgVbxiH9+2lVQTFLZ1JNGw+57LTPgch
YlPRD90Jbsr6J5rgKgSM2OtcRaj5HeXLeGfYvcZSii26BEUbQ0vV27IowXxouPDi
wBSFlMwm0Zy+leeymJc+mDA0u43D9ishH9IE2SnZuKu2fb0ZdX4a4+eCkAQQnyfi
MPgNnAT+8a1IS+zfeaT4FKqsb8V69ovRZKfCen0wCRnEY824ClglfcrZo8aEB97a
FNTse1RlbDpAtKl2P7Ori9AN38/BrW2VuVdxNGypwNakM/PIgkChu5CmNnPtI8Ov
iG+LaieBvAC+BUS3U4WrI8RzqUpRlndeS0dCp/i4WonythVToE5nRnTJZtg7cxbW
UcL9JnTNoUSBAE7zZM4/pkSOxDkGMIxhdkbruCMLHpRue+MuXk8fjAkxyQz3DM4b
qxR6P9AYT6KxX2qepW4lMlUu1ZfXbyj/jC50YSec9ZrOzTmtFYtFhPJPHhLKL1z0
lAM1XKFlE0mS1s+P2WtaO8v/9JZKFNA9w7TnvdG/Vae3IrVggM2sPM4GgZHwT9O2
m2uF/8nF/EUOym9LwejtcyOQzXVNctQXPSYDrlJKxPVH+QScNAEKJmEt8/rNUhCI
Be2EXHww5ggeKVOqia8iqWyGyhftAlS2IB/HaqTpJz1CAiGMmHNBSZ8hBiIfsycf
xe4XgzfjFyBeuy7DK5iOCO+Gmq+kM0tyH801HIhy8r7bawn9szQuXruh4YGfYlfE
1GdT3cnindapLvpXbDeGBoqHdWsIMyUt3q4FVKfAVyOx8PX855jPDV1YEx8n2Sre
HTXiDsYQKicqauptZCf8414Q3445Oi2usWutcEAoGk5YgCs+8mUEp/zJs3eodUNN
BWvohIugxKPqVVyxbhqDVZSt9tNjEc5cIOLi1E1+2WENzo0/Y4dg+zRqPxE4ALz6
gKUVrIzEo7Qp8RxT1JbP8XrxsH3VpU+NZ4SbO40ldle8//xOb3TXHV2S2xkAtR59
DSum3M9OrPzGyuOYlhucrEgSEzsUqeRS6L+AYmhGanPD12PvdC+cuzbaqW2JIEHp
NpPHDZSpMB0+sfpfsPIXKCOi8omZ02NMzYxpEQ1LaXB8Y+P8FN1JaB/ItZLV7wv2
4MG+NDh9gxHSKGtzNLPZ5CinIZRT8jvTR8DamsN5lH4GrbHjZhQuKn2a1benoFt+
sfZS9uI3sCi1Ry1Siiu5UhtHadZVyI92BeXmnoU+82eoByGcKsry4HmgEQzvV+gw
QZWT0CN12W6TfSrO5qBp6UMkTvO8XgB4y9PkeEjUbK4zXXbg4BAXzPEUYi9khwF9
o0ErUOcol1tFs8+/gAmD7zbwslqNoDGGt7pJw5IYOZBtZPnSIqMSgdF6MAyWvVD2
wA5zniy1v/iZa2GF+dH2neQHA0gGsgosCUwI4ONXocIAP9+b5KYOQUU6c1E+Xy5o
iEchVfV4koYv42CE9TWaRG2/n8BaOAazWiboPrLKZbQutWU408BuGpVOU6Z3r+ER
4DPWb1u+P0F6IV33RQS4kgkHT4bFBpjmHsdw2dottu2yuLOg33vR7lcS+rlrAiSt
phns9R9GqS0hKCGaVcU+rhkwwDVI80iQd6xiH6Vw6ZMc8rz5eoP25Q8CxaGvlBVN
yJPF4C5XYPogRSJ7lnj1UMi/9GSZfrn6P0G7JhR7dGqH4aOe1mgNDTBO4DJS6Dcn
UWXplEt1uxzSGiajofmLLgoRpQl4wNvNgytA8aVuL1ef9F19d13ONijhC35lDkCv
/xqNF8E09IIBwub3Q/jO8ecQHfHYduVy6Dns2eWR/gDcp8eEz4GGMhmgntFyWsMD
nJZXealJ01yIbbaDLz8GK9Sv1hGB/om4GCFBezZ60nxeRpIHBQ+B8Zd3Na96JuVj
zUaUfcjJxweoF9D4IxGHeejnn9HOf9PkvpGSfI8zIIWzr0IKQZDuE35hBvEPXTRC
YOeQpf85lJ2Zs/3vd32qwKzb502ux5cRy00cfFzsM+AkAS/SDurvLxJf38ckvuSE
2AvXnGzOYKmTlxrm6gkgFTJrxN1TZnHC4g2zcTsOB6wcPUq2+qKJFDqeM0Y9r9vT
EWfOKOVpdELaC8/j0nJRVa3bxYEAuERhJcpsGqFajZuF/Xi8T1Jb7l0o4UMNSAwJ
jSKSIM7iASsbuxRq4PnI6qKNvnj1ZYPS+h7Z7aJZm7VL+ouzq7758Jv2Cw4HfPxj
Eb6C6HUJKbS8a4Ma6PUoTyZwLLg/CITrB16rqdwx5D4taHfFTbmrTPIQtl9Yxml4
dzj4p0frLoc/BkkT1/LB2YZueARsz5fR/CyjXBesBmUuvWrPuImo/WYxhXlQePzx
xNpC+xgLRL4/WkZpowIklswKfgzP4qJoDFJmP1vxFjF5SI8RMXEh3gg7dz5aGDgh
sDoEWbSA75sxQcZlHICfoJuBvAJ3JZnxlvmYZXzvnieS/6HtCsfyqHRGxjFTPwMG
KUN9CJfy6Yd2tPJCBsu/bfXXHu7EET8hA8i/DnJGho8OJNIJHtFtRDxfFkExCDrI
+VPAeG/aIzT81q5zGIuDvgdaSIFoZjl5gqMuYLx2FQz73Gww0hIljlwByJhxJxPD
8u2nC+3xSvGFsUwkkNl8bzEJdrfImQu0QvZuZDHw4c3lF1tDJej+k2/5b5kEZ0Vr
1VVUqtZc5JTmy7VLoq8nm0DzY6Iw9nr+DTQlbCVdCuUZ7Ysi3a155K6H7+Nxo0gN
xXbYQnhmQUMxFGizOZ/6YXKARM7ZA/c15ljUtm3YSWowgI63nmnmi8FlKFKNOCr4
fzk+wyj/Mc4u5ezpT9dM426O6cFwhR0TEyzMoKiLo3xTthHBAiL/ROf5d07ul2On
mKuHFQjCdk1KXrz1qugWZdq2hxukrCw7ApNg4K6R6+j99k5hdD8dW1bndPZecxKk
ytxy0HTNkRI4dV3kaK16XGuDwNrqhCtgDmvX3sBJsZDEQk7gQy5/aZvH7F68YEFb
m67lNoCz3R4Zkki2vhRx2o1TcJaYClaVqHi1RZWSM5kFZLSUzOz2OgM1lKkdTpMM
WhJG/z4dbDqoOvkCXKnaKSSC5CmtcOz9KwZpzPQV0fx9kkSyO85IeYDHoW4W1tvB
PK75dFNkit1bFl9DwRjYIhN/9pfiHRmomIntozVVDA0Nk4nBcBlif4QA7lIbIMIn
F9c0N6FimJW+YFXZLrSVxES0U9pZxEgVNLqx5hxEZqd0y2HAXN4vaQc2zVU5uk7c
0CnCFjZT5I5cM/pm7Gm6xepOzGP7r7eXRvYtqJnhMjzWBYENIyOAZ1cEr6kAwMWL
fHSL2H4JiftGGKbc1TRxYokwJK0sR9252DZAX0CVAD/4pYTjNUB637fFB0Us9Rfa
Z4DhTHAqpa3+OrMps16rK3/6RfPgPAFUJtm0umzy4bW3otjeUEwvwDcGrAISa/dP
Gb7u0x1LI6w3zszGEyl26aBbHmej1o/E5+zUyiDWwmamA31shZFjK/GwPgsAvGzJ
cHx8AR5Mk0Z8Y9OtLgxLv0hogVidmltJrFBewQmjIj1emPef+36hdLpHjfFHufI/
T1r3lVqVWx6gPGyMVfPmrwewelEMl4V6UAsEvzsmx9YZR+URkl4g5HHec7sOQ2mO
MvFkNPWwOAHPHj4/7uRed8/2SLeYzZjKbISfDGOVDz5G1FAEKmou3bS7HEgiDo/t
oie0Wz0Ox8+xAOCZJBIYGFI2rV6AkUvkH9w0UOHbC+LviOPi3ky7SG9HoJA6R/Ot
qebHocrLI7EkohkwbgnhxdTf0vaZXv+jI8XlHPLdEFYIWrUrSYZqM6FyCeKTH0Hd
tTpQ5LChaimEigExD5ut9wQrtpQt6aUggZ4KFUyZ+lRPO3QONoS3wQtUtKazBcGm
2yO2cWjY3cetebzO8pAfSW7IxJL1gLuMuSfigeK/nXeOWsYmZ/u8uUVLdiX53BoG
dH7scPnM9mkcblPJqev06jWFbXM1+YHX7+LkFcxd9QXOINFUBffPvWNr8KZwwHHx
RqGp93+0rsq/vsO8mbDEP+G4v/E6htaOO/BM2TnrsuUug9Xf3zLjFgRqt2ceQyVn
KvGu/6Y0btomcCzfs8tYxmVnpTDTAqk3N48gUQodxQ424Za9gmJrl9OYVQO0CY/j
KIpRhgfB+e4XjIACmjGCGZywIG1frSGZqgY/oCsTJozmc0MEOa4g6qFOm97GbCp2
wf8u8qbyx2gzdvzz8t+iWl2DUiZjxYY7NO7SapKxRjQvqp4NTVn83Oqz6TdY4wJQ
IIxaYes4B7VObVfIAEH3R0NANVqNo2pQAYWeezTonewPEdFdmqxFSu4y0sUbj6Ga
sSexI0P+kJZ3WjcL0JImc85mKMrJZEpDbjGYRYU+r4dAXfEhkUAFlfcWJ1dOpLhZ
YLSJkgKVasCsruWo75/OngoZUnMTnBZ2IYJh3vO3V0Fh6zD3GiVmyu/949fQ+MZF
v4lhTWsDDFI+YE0028T5HmQ/YT7xGckEJs0KvwtseVgmKNM7JR84TEsIfKzgz6tk
PO9wx+YwzaRzz+v70TXBouQDIq5T3cFy2yM2zSk0QyjldbmmKbgWAGC3RolzMSMi
HFJZz0cmdADCFLDF2TkgElzkGImdZc+wIsooQbZemOZ22BHvB3ZUs6KcJfdcYcdk
P9yiTCchfsB2HVbDRusaVkx1BGNt65P080ykw6zL6fFmOICgYxBVWWWtfXhxq7vV
YffLajF0bUA6pkfVKsCUQtlYAFPXaZhT94CpdS/1d455VxVFuionbLwqQMUe/zlF
+aNuEhvl1rBIX1e82lawQ9H8Z7lexHt6s//FQBwTjcYpwlYltFI7yRhc44UV3ZTq
ejYbs7BKhlpP3lBFUgCbOeDK1Dm+gYPodTf05Qk8gIQycew3zCfvql7wP43/zjqL
x9TWO54CHZkV7nGsiHFTKPCDz+h8wd0UsqmvqVe2YG1cYQT03RdgfxDxhTV74BpN
MWCKxs5dYInRzPVcvkHaGswWuSlcpp3wtdMRYoprdzEA7ImZ4EINBuoZrcUtenY4
yaGYmYomrsI5idxrbCPqI8p2yb7s0HJ/kPSpvGL/FKvtKnWVo5laqV7/RZNqSowd
nLKH0x9jyRK7RsL0+fVOyWI73AQubXnA6ntKPSlU0ZV+9jnutNkXHkkuE4mZctr5
Weq+/8F5EKePOZhWV9rcWlsBxRMDs/nPXozvy/yUcySSaywaNHtlgQUGvt3suCvR
bgwAuu5x6wp9LSOsXf5zI/Jv6QzEVIV8XgbotHPMjbHR4/JN4jDOjsfycOFZ4Kq0
uCV4/gfPznw0XVsS4+JsAsqB6ezYhiehRirQQLTCxtaGb//yJXbIveyEF/GHof9Y
UOfXk32KBYLi4lwFhc9L9hAhpypQcoH8ylHwiv+dOLg7svdZIhAw5HUGfjh0e2YJ
32oyn47IG/WA4F7y6Z7L3wEkLGSQmkIEPiaXsYAnjj82WDX1j/GHKN0qN8T1a5YG
7QL1uQCM8MSYphByU8k9QSfzaERGoPYtTcMSY80b766fBKrInKEiKb5r9u22ZqmB
8t/zOduVkFiNyh5N7aciLqCKF57L64BD6m/uyG4Kf0LW72Ciu00T9h1zPOKKAN/Y
boMLOAyRJ/esq/2oH6gWs2W7hOcNbBGs0TNuZWxF+WeTEoocXLEEC4cKUKBIWHsW
wfEdKmr29zqVsUKPdB7LZemVRTulWgaaICBG5uI9uxAMhuvxEnNssrI5YjrMl5oe
4J1IEAeg4Biaa+OCGMxQUfeUSjDInR4OG/4aeJnesLUocPaqjPrxiOTa7K3NQK7P
5hHmKHhpVoy5esB2oStMvd27G65TOCD0Tf2rAmfW1v66s53Mlzkv5TRlwxcmqjIk
dbobH3A+U0U/zP5+ZLoEEOVBqof1qvIJRYyZeMliZiF7wfNKKJmAR9H28wMoBAx0
gP5LYy6LpuCnVCUEVcAdQnWesb0/7S+LLY5ldOIuOygY6sZNLPWXY+58ntsNyzj/
3/WfHvfqwqebNnYIX4AM1yPcTH63aEuLdjLlr0uKLf76SIsE5stp85ccuW1qy6pd
AqHCcVgs3OBX8fF3G3LUm6mxtHJ+kn65T/wh9gnkbXIhNBcAYklEq9FWEtx9h8vc
e3OQR50VDMVCa2eY+we0nzxg0jH52I74+/mkVFQyD/t4FLZzuk0Ss7R30S5e3QT/
kk1dUT5ZgYrOgPXNGsuvZi6EQb/5MPR10HLGPj2tSHcRd0C2adzJFsuwHTDTOta1
qMZoGFDJkr82wJ3JilRMsU53w65C4rUBi9jQIFgNStc1Dpz+WE0WxscTxjZ/wzO+
L5pILWICed2MwN3VeRb9X6Wq6lmFhN5rsDrJEDapswo3EXuxUxMFYKSXUEYvxK72
Si1qAd8p/k36hfdtWRWo5okysNfUDWeeZRv9qT9rVQidIHPp9MKWAwjbxZQUPyVC
cweh4t5hXq+sCaSnPHRlb0X4d332PhZlYMxK7ZXPTIRu5H7+fbJY2Z4XBaw0hcoR
r+NeGzNIcGTAuwKujLAIgv7gxn4wrOnKduNH8pj9Gkpu4eHorDWDFF3vRbWWN18J
JmXQ0Ol0gS49s2ZnjhJxtkVPrfp9LkTRC0qpKrPkwClY+oqdJcN2xUZDnaCy2gzj
t1iZS5sBPLNsD1Q/MshVlxjPATd9I7cbQjj6y9gZOW3Ki011uLIbchQUbRu1bKFH
TUBYNt92dH0pZbN3czbEpkVVuj6ErcXWUpQ8W/XWdJwtoLdPKii8678zoSp2+CvG
uXZpHIoXptjxGPb/v8nEBzfH27Jj6cOuu+/8NbagcPmWSoQJxKtQ4NdZOckxJgam
bAOVBC0EdbMk2hTZgmQtRFAHTJObpFbCAMoaqBOOKrVSGzTfV7jtRLj1CGjYtOir
aiLzcCk6vi3zs0ZLjElZzZBjaaz2BHmOmfmiyk+r9QV8ZGTK6N5fVfM4Kx9lri6z
oR/DQAouJx8qNXBTq9C8jw1X4BAUxXEs1kx2AN+/i6WaM+yS/d70Fi1YPqc0O+V8
cvTUnxSpR4qheVMOe/M2EuUFekpUdNoGzij6GSx4L7xWnNM/lZacLu8VNunFuOI+
T+10qRxgHDhYIJnB0l4v26CpnFfp365npj+CLOJqtt0dHKQyv2+lgQHy7fJfog+l
1HTOzRiPn597HeLKpH38uDmrc8lJk1nsR5J+aCqIKQ7EdfWVxwIF4P/uPsdoQPK/
NSoFLc1XsnppfAt+Nv5zALeWWoSQ2l6xFR3aTDTFut+9lDNnrVeF1SpKrTVfz6eV
gkH4mlZNloCu5Gbt6voDs0cTh+RaUq18qtU4ULVOQkoNi9PaX51nyUzx/ILLeJLn
cHfiUjHwKNpe2ICtzgqkiUA01FPWNVoNwQErW6ZEcpLadETy6GWiwV84Q23BP4LQ
3jXyTW09USPKQUX73rm3fbtc+1urDuf8KOV8LtchovBlF2TYja3PbLn+l0mwHCqd
dnt2vBvCx8N3TvK6oq1dUvphUnLG/IK1WPHlD2MRF/0OzVFYFQCZa7P+TmYwOOaS
FwXlfeKnYOSAGp99N4+oP1C6qgJhnslq1dTE993NT+19lcMIOaMdZXPHyK6syPBG
rYVOi5jMgayTt/Lx5qsoBhr2wMDeyScAq8nmPd4d6tH2lNJDHPIKt9LOzT8+Wa+Z
Y15XtVrJ94nmCARXuQ7LsgSWwMZ1bueFnjTiffJ+1iGZpLn25gLUvxQc+tG4vu8I
09g8lCMa/s4RRWuizJxXV91cYSMb9MhVjTCegAW6mrsNjPSJ8s9tKyii5Yz1hcSk
O3ZVw753eW0mKaQR0gX1qtpoP1BWDlx69+D/zIFW4ApJC53DI5WXEeBLZSsHAAoA
0JMbtf+PHn+KV+JGGApCtyxifXj9DYNs4xy65REWX3YrG9qEEluGR7qzLSLCUkeH
Y7BkdQiCUvAoWZgHwN7kGovu0Kc0NAPClQbqp84msTsUIhWXnQNKIjVzpJJq/eV9
3SQGJ2Md98I5GOEx9rVUaqjyc8YOQ42qf7WRNdKK8qqsuijaE6lbIovmqDj5wkyh
ljeWX6wZ7xz6IE2yyv1IXZKtVrdTfTFsLCo0nKL0Z5ufNcFTXV/rj93gEStPu75w
5XbTWwLn60owiNPKQ+ziSGQ5l5iY9EL1Vlcj89uNahTI4VmSX/gmPVJ2lvjLo1Qz
mC5Yx8BBBR9PB3gcHBNXfuQQkwFUT9xaA259sy37hcqdzNL2eZnWz2ml6oyrfCet
OI2qZgGx7JEb7caRD4l4X5tHq26fN/RSp1iPWYrwmYYBi7OT4KuJcEG5sN7a7LMw
43XTGnwt7atbiguFn1I2WnMDj0jlCcUBxSfOVkm3a313achFVg9jol/0s0cptZAo
j1S2gCvyBoKBcsgQTz+dTg3Z7DFCWiGRNM3JAZAzUpWwzaxrzb6GAVj6XaDJv4V3
4t5viPk6QwnVCzfn6gnpH81AHX8/rSkXtc2V7bIF1DiL1PxW1oWelvL43r/f/maa
4ofv4VFBMJQ1m57va4u1ZmOn05LJbuPo1hhNvQxndjAp+ZqepJ+L6Xs+XEhvvrDo
Jh3N/Ksg+4YvZ2npt6AtgAW1rvNeuFENNyo3f2ftVCUPvyEB2Ba0VnnFzY09/YTf
elRN75ShUz71U0J8egif9Rk/66oG02mK0iQDQbCN4i1SIJ0JvSK6eKqyOZQm8BEB
GQ2SFLTFGMIgfEDheKzhky07LaKaTPavYiuNRDFm4Zq1pRBqJgCxINQAoR65COh3
iEpvzVMA7EmDS17fXe+D62bAaw1gpiyXEju068iusK9jwoPu0YJJ7cHtAOgCT/oS
BEqOltOHP+L6lmEx17EpciAu8Upks7UF2S14xFEh4MEUJXolH5/5MOGKOrUlHjWn
fhSkM63IVn6YGqKnzZ9MnuQBz0DqojcssqUULpjy4R5UEw+90r5jkAmUADGa6e0f
oJplZSBgMCImWY/+YuJS6cfX/tyhcyAyimMoVPO2UDU5Uqen8ykMuQ+BB+P9BxgJ
j6q/tY+q+AdyfGCSnEKFLbA2GsHcQhovpnKb4NyYU4yGasf4WbMExosOyfa4GFFm
QV/hl2v0Jm3P0lHNAFucQvCUQLzXu7WtgmNvcCRfRNr59bauZkzUNKqgI4VzDShV
f8zU9Px2AnP35NyEq2yVxxZkoeZCQWNhje1sWxNMSPkn0MC8aTUuAl9ktwsiycV5
YBAj2ea7rkynA/Q4yewiQSaWCO0SmOd6R8wk/LNV6sctpJsGsk5VdRN3PY9UD1Qn
cc6cVLPPO52qPaPcUaBwgZU0e1KBcuVzG9ESAuBNXfkNxIvO7wa676bWpaWNct3N
4qrheoQ4EmMPgasjOQVGw6gbKn0eVRfbbEBXr9RI+kMQHFfusjt6cxjdhUReA7N7
O0Q6b8UtMF4MRzranIYeGK6rsxxTfeE2m/580w/IWqSw9aK2idKlVBEoL5V9WrfW
T7ADPnGcDHPsxbMjB+hK9mFIbhrIXXaDi5MmsKt9H4LKEZvpmeT1kp5AMKKOOo7y
73eXVVy39kWlTuBlN7J5W1ZozqY3czhaoljmY8iPmINFcJNPo56mxdiXSK98rY1+
ed+okehVoK7MrzgCu0dF4RC9dDsgvLcMwmah6NsaQbB13fO4YQTKf5WLYOMCSTMO
P0QUmbpm0Hq+O1eoexA274RS5orbz+/vgo1z2vj9zBJSkxn9WQoIArrVNOKz1uu9
eGKGMA7oIrRya0nrgdefgn5KJO+Mk1LNBgTWcDuc5ICHF5PgJTK4+g0VBRUvjEV7
IybaeJLcDlvkAb2uIhI6WP8BRza6Pw89X3ACw4lDO1H8nSj7gC2rJ4H0PWbjlGtQ
Ry9Jpl5A/T6roDW0dnMSRc1QIheZPvoMJ2GEZyCare/n8EC4wKunNngbzj0FJdyg
l+P60kUNLaxZIWiTqxJ9LZLTJYaS5vUvuFDpxk+Ch0ICcMa9c97DugjVL9rCnwbh
W7AyICkuAy3vhJ6FiuH+XCu2dZsZ2/v1yYIw//VNCg8cnPTiwQnhi8jTWwRS9ke5
9kyj6dwcYxVeuuLt/x8CUqiBJe29+Nau4r2pOmiJzaxAseYbzyfTzQ0WbKA8UM5t
3061mIjOr62NA0hTuy8fCR25s5V87AXnKqCmPSQtoT9R/rbCcnV8X4ERKoN8DiIK
m3e6d0+c44fjESk7lvebLhXYIFFeItz/wMFSyMjTQBarxeetmDzD7wwew4gASrHg
H/lqs0iB94JYRFVVwnsmh7QKuunFKFJ4FcMeq5qJB3J+SslnnKuyBIntoxx4oL8r
B28+4d9CgKpudKEFwJEp/KYyE+dWgAbKRaNqUF14K8LQsQuQdFFZrsiPlSkfF5nZ
O7l6fRUpR3KyH+qFOUFASUDzuWqCD5GukevOMWHvtDQHKLW2vx0lcNGEFhaw3XXH
mBEPefb4rX318AschuqKw9POWRCdYYiCNQ47goOPO+hklT27K9ThwsxiCBegDJ5V
6HR54iaEEb6IRBLCetj8ntN7QkWjLf8UTSokwlrS8EOHghkLjIeMD3hM/CnbBY8Y
6ajQ7wC1zI+JM4HHF02KBNxzPUBWG1y4SKfVDD5CAsyt1NQDYR865/9ua923f3ap
1GmMZ/W9rrxSUOIOWEjbKFHP0u4bnJupYt0Mly6Qp+9U2fOBgbB2Nqp0XIRhtO+Q
TuIwYuxOYKuuOC0q6HAacccSk4BNMGqoqTCBSaPAU+hfeWOhXJVi5DJMoBRy+HVs
PsBieD7DxcDSmYxZgu6WQNsj0Ps6N3KiXxXRdpzrfsMpKbfTZGzYvcfFVd3RigPO
IrQ4ygJ65nWhvfEEF7gB316RxKmNQBPEy/L1QVI4Uj/MPKLKQeQYwjDN3QbFUY9t
EPep8s0IUcfyS/jXkyq3C/q0PVJb6jW9m31NKsscYN/KCIpDK1U4+jUXK9/CaPzU
9DfjfBHipJghCYplpHiTrRZGwPp6vLlozvYQdLYmbPC2zVUUPMP6eR9ipUjdOnA4
pD/inMxcTz2EpYu9qGaj0S/XhL2SSdb943R36/W8YeY6+pRhwCj1jtI731DfS16q
r5BdpqOgH1phsCaardbW37NqstMoeYjURBEj37nK6nAR7QmsNjvAEiFQQ86wTrYE
G3DqsR7Aiz+EXacHIrmOqwXPElajqxd4HtRs341Oz+B/oXp3LFePRf+6G7xFHSWJ
/YjJkjhoYbgfbJu14QIuG6BZrIs1FhArM5LTd6l8U8x8ZSHERc+dHOsdNwhU3+yH
TuGBIoXE1AOCPZFyGKIpP+I/z/UG6K+UsPJZ8oyL3mb3AL8+zyMlrSj4OWq010Pj
6Oh2XKQ12DLMXUs15G2noxke2ZgBUccBbNpCK5sYMBwttAgwb2lgCODUt5OGXBQM
+fY1N8xG4LYFHz8jaFyEPlbJ0G3w9J+o8+SVeckJuQ2y6NZCeeZZ4bhVCiq8kxvY
/IbakJTaJFGDqv4rSjkEZYdw4u2dkMZJ8oWgLT1LdxptSZ2v0NQOBgIc6BLCtZLm
w06vOuvE/RKeDIvR4b3uGg8lKU+IHG2h/c7GyXkYok7J9ur1vvj5CE0aM9+nEIET
1lc3ECXlEU/BsKozD8lfn8QnqqKHttE1S89xneMYNn/9Pz5ezq+R1Wei/1l/p9Za
BLMSDglyESiw8hU2gra6uW/b6YhW5ifkrJl0ocHoCy7s/5lgVMqrjXaEtw+DYa3B
B3cVd3GQsmxbzNgqXeudouXydmYAyuRdDfNTEKTrwBC3h5TrDkk4Px023I0S1H81
tZktybnJi6zdyOMtSuzTFt1gnRdieVlk1ccwrGGNXSOf8h+y+4+9zR1PeyMP7W0N
pT894rErLuC5/bFiXmuTzNTNuC3/fFCFStoD9/KH+LkoP1/8+KT6uz3LFHTwwhR1
RL7YzflhEg+Ul50fNGj7vyt9OsZsVsJFGjWdgoGfJUMTTNo7DJNi19q5Ubnw8/tA
Mid5N+9REwLPfAEvNy5I0xfV48hH3K40ZVsBdEfIIHKb0ndvY3UrPVxVB7ZrI1hk
70KJQJS50kv3/hxNgYUu1VNLFmtTxQYgMLfprizX6DQwSp/+3lxIJ+VsmEM+w1cU
SR1KkjXsgMkcm0A5+cfNfIC8nZUSMxKZOziymj4GVntP3U8uXBuzYkcABRLuJhDr
7arYExBY08k+k3jDVzdS1Tq6dD0fmJCo+cVCvgB2zezwWpCwdRaA12x95OcB2Iar
yj+kYV040Dev0Z/lZ9xIXcSYVMNcXrCzAsmraQSBLzQsOoMoAMvZ6F45ExGV4ORk
LBBEgaHBoIBv+OYbJAfse6hvFIK8rkQqmGZWRTj7bxHV4/AymgCoKFVasWHE7EeF
D4SZkp/SI0/nUD8J2d0nrzpusTKs6J7pjP+yOSUqO80AyXA62KqfCvY4FAy35ef0
Q3nPZnlu1xW6dAPZ5BWFpEjk/+mHgf9n2wXnCKmHxj//SPFy9i3lTxNdj63rlCUu
ZWUNRs5rzn+CF/1i+qbq5xaemSTE5uPAaBRdAA8lSYB4nKkIoRqeOvpLOffbrIi1
+f2b4WlKlykHhBu7KOa1qk+rJgFWgU1w3Wt2uU9R+4SVh1CBbZ8Ry2mIcn2tioSQ
s8jiSJGJyPCxuuyYsKzWfW/AfpFHL4H7VWOzdvpNVyORxZwbDoDKqvY3bq+XC8cf
uusrfXH59prRGXcCibZ0OW1FmYR44zu9pg9DotIrGUzpnqjVO4QejI8AZAhPGjZM
fgZSqEp143/snNmwTSJTXd5p6tZ1ip7F2wJm9KToSSWs/cTelCg3lPrS3QnPPiwx
T47Jz5C5ECA4yxoNQhpTaoTyur7l5ZvjdPjp7MKqezyT45gK2OWBgQcQTeNVXMw1
oSAlWw3G5up5AtQpJfqOgBSWi9V2JkUQaCIc9454NXy6Ora+1SRY4GDAVsqAcuKW
0+YYyOHNrdDcXRDG+WJk83Iojyu+sG5lUc/7zuKV9XpUReUlRy60/ydYoaeJUEoh
Sgtu8pTmcSyA6LPSPp7ieRp3une/WE0we2hQf0HtbuDIXj3Oz7lVxghua5lH1Z0w
NindWyhQa4Ljta58sB0Z+TbIGl/IycacLPfJOYMi8a1eOuc0zC5YfgLJg5E8RFi4
anRRMFbHag1f6chJzJVvl/JUEM4Lo6kEx/Hr5mBUG2Wvt++j2p8cjoobQu16ylv+
QR7dxrkLSwzSq8OO19ZvOiss9uxCM1IEFcIYquSENa+HCRHSFQGfgyH+rFdY1Mza
XJ73zVFjYq2Z818Eeq+nHfeU9EYwwzn6jx8Fg9Xz9ofQQqbtewtzJ1qbjajE0FSy
CZT9WXMmvwQ69iwIlLMzjk0pyYwrbclWTk1ZvlTnUSgNfxRRNF26BhdPBo3WsT8L
z9FUNS0mGQpi/AHBXffCVTQB1BCc4pi4lLbb6bsQNTLovkvNwXwOQKNVLfq2GwsU
rVfmBwwUJ/MnVLC2Gh63Ukk2K+EvJ/MPY1IMLCos5Yh8h3EtzUw6qqc5pO2Rg9UN
hvUPSj0gnwL+2Vw6/Mh+1FubsN5XMGU8o1keOfx/uukeWg6pijafFKZ/7qd+/PM4
+Ckeiec1fvhJKdqoT50hK3XW94Co0Gjp/VNsmcGDZaGataKuQPFlUXpl7rdR/BrP
44ykt13tSQTOCuklzvI8BLh3f2agmHpcNmO3H8B5LbDpYnJMkj3988WKCxQBQZov
EzJzoA+QweWcMJs+jBaVzk8usoot7WbAHClVxuP5H6EhMEWxoN/N5pRmYr1K02xb
2YLeO4YEQF2SuvrPCp1+3w8f8cH9dfa5mb48aUYBYP/AcVzoak1zMe9Q3f8Si7P/
sYmEc0N9wE/GmtWjbLvHmx2h0OYB3gwasMhtMHBzu4LGRnj7EujxgV33njH9ABfY
IMwwM9hmFKIcDjUGDceSapkc9LKDAI9YHhQPX9e6xADEoW2VuY5dBH/BTD9zayPP
/6YusuRVTiDvy8IN0GBzu5fFE+OSFzm3rp9rT1BjDZz/IrWO+8iptTO9C4viEvv4
TVElG6Om2RvwOXDNcd+qq4OwrsBP4h/nO40Xg+EUoqPi9Ania+Fb0u3ha0tXHGla
mwz1w6H2QYvviPsMUbuFCLg7e++Z6V5aJWUWmhvw5EzNS6zWGZD0Otx8eB167XDp
jtq3a3NaAMbADCjpSeaBCY4hM8wOluLIett694U8VcbBmHGtOK65CNfhynXJcfEz
Kl0CfqJxG3odpnhFScvXSDOmoeFrGkisiO1PwC/N+PU9RHf8+wtl1vagzukkzrYd
XNMkpUPNACAgXTbbq+TdARsgck7FdKn9LjE4PbWs+rWITbY1VFUSCU7FuYvW71Rs
FhMpj07XH2MmAgQiYQAaJReJlnZtUWfkABlTj/8OQ12fAOBZ8telBlHr1uIjRKrA
9dADQRCLzpK86MuDHem5RabGay6MF5zezeTweLQHhZmpj3D33crSGRDv5pBSQWRk
o+s8DhRSfOboB+0a8ilBea+RVOD4o+bPVNzl3wsrUSh/WhSAu4NJ19iLGG3Y93Qo
KEbH5fjrlM6B6OofO5JIYcTj53l3soZWswU571RsrzuTAjrq5P63boJ/z7dneec8
TVttpxtU5sEDJF6Kgpwd+s1rC386kb68tTSLuGwc2GPdg04C//dbwzgOZdgSC8rq
ogErKcp3EEI3Ak5Gz9szA2Zp+gicQ5wZAtoFKH2XJdP2iSprDMd6kW/uV0JuB+hz
Hx5LWXPQb/kK6eFdI5qTPEunXDnoyAGJjxbpRhw/Y4fhjDcbyt+5VTOFU6Jx/P3J
dRCMGr1xB7G87p3pOmQe7BDQAT2KjGjOrdcN4D04FUrNtoop6DZpkKTChy9Mq/Xu
KrrS7k7WxxMEexPX7lz4a80mcNlVTgpO5+Ju20SMjTpnIw2WAJb7QW3rjDcJsy1T
zf2YCgUP7EdqCFsjIyYioj4Q5vEoM7btZpkfQaAEZMLZNebbRScEiasWxCTpYZPK
OemPkNKCqK42GAH7CWVQyMqr7djUHyPIaWpoViHPLGGQSdTlPNnhjzgkAGrLVC6f
00Io9vzr4pcNF3ftijTBvMvEoP4r7nnqkRmX2/3pWRxMkAMnRWGilYRIEdmdyRLa
SMKfGT0FC+S5icUh8xJ+odoQddeoUcGw6VCCX0NxNbL56+fdp8dFu4+j4+u1stYZ
uDUQpOlK8ErbfPYpGOXxiyjbBRxH9n7RCOMjE3TDN5OLAQaxHxtI3/Xv9g4G493U
AVu0z6bNAHmWXNcfhRjFveUTZJth4f58EwWou+OkaxyJg6c1vTDpKhieW7Y3Mbzt
dAlmzICMOcJwq6SCPLi5bh4RzAUHTX0NENwD4n1srCbCoC1YXffFQyWhTM0faQWY
EAS+CsO8iigkE1jL6D+9+GnNTYpXwMfdNc335OdeWY71RUvlz77JquQaeff8sPnb
2/IEcyzYsR+j7qJo5L7CQUtYqPCSOdeLE/TF0RIpZ+ktPGai1tPvdjd7uAbLNB3o
MQcl53559u9oDSegKlzM0t3HrITP5ZPueOeO+zV6pzHUvC7tcq+bSWE3lcmL0xo+
Dq9ODkQa/nvDY3pVCsrVWabXYs4jviO3ficuhpQD0gVVUMqjn8uIkBshY6oScu04
MHP7KsYd6Yf17yQJXBxcto/eNoNbAgWBNoDpVx7MHgUFYrYGjQo1J1XaO2TnJN3/
PxJXAr5r26IRNhKVnnWd1kHx9RFBKDhYU6z2MtrEG9oMImbqkUjIDu91hfZMyjcS
k0MaJBf72WlxAxeqDgVikyB6849vGtnz+ULEVY4RpBXI0rTsbTvKJboo/6ovAWgi
8S3ITPMUNxNkYR1P2M8dMHPLk9M9scy1CDe4rRZFW11ZZoQJn6GvYdQIF1AD3/qA
GRSoLbBdWGSbVYEX4R7BSZ8oz/lvhztpeLubrxQm6NR5IvExfvzLucw+RtYU6i78
agpEC3/jAN/v68y335C+5Fn8+mBgn8hzhdwb7HbzBIBOnpp1iJHyMj3aC8x2eNrv
83supLNyj9RM5O7riuKH9BBAY2QjYivFdORxDoyWgJ0cA7kpa3qjpK33qwmTQk9n
B1bAqTNkFMRPHrmkSgpWwdYgfWlNxFwpemlUOi9qDDfHnA+JZvfJnnI7De7Ar0z4
mFpJwPcKzT2RXkNWAZLl0dfpDXYfr0IvnPQBQy8TNOsVmA4bdJ3/VIBryybDTfEj
ChVDFzM1PyqMwKH3JmV8Pqa6Vruo9T/BYch7+BfGAM0oNjmGyPznfiIL3VWBnRny
IHp13pFEyxtS8OWaN4EPdbknQfU8p7AFiMt3/G79S9slUM4zvtWx83n8UPqisWj0
vvfAghiZOtwZZMk3VWsLOIvPB1RtV+/jR2Vp5ojchX2SVQRoD9+zI+z1TGZNDv3v
FViQyerOVANGZ7qrb0Zxz/4T0+pNJPRVziAVMz1XN0DmaGUp7Gy7TcAOpbBtwXf1
iZSnHOB/jjmAbnr56jsidBItTvxYKJ2RB4ZYSPZwLEl4y//T8qXjbq8rmPevKOHY
UyPq1ua7iLoymEPEysw+asGgSFGXuTlABe1O8w1Rg2blnR65agoBHYPCjJHN6fHR
D2dMK69yQ49C1E7omj5BxLgEqBnUoNTuWowaYX4dh5D5wN3ySyYIwVqQ/P2CvSjG
kmr2ftBemOX9S3C0UGIyMJsVoa8DYj70qWGcsNsc5QsdYZertBOWIAvv/j1WfPSb
uXuMLdHJxrIYFYSRc8jDme/b3FN3VWv6mM5PwKaAMXVZHv82DkCzf+DSE0JoDO05
HnSWY4SusbSQgG8ifpw3T1sPDCAiX8DzydgTfAPH7ASEtLfQhP2r2n7VYX6oYp+1
mvRwqf6LteKNpLY85/VjG5aaLfgNZBseA1hefBVnyF1WVDAHSr3HwXnhvcRvrlfn
CWVk8V7HSYitqnnM8jd5xHZPf1dxm03o5iCXXmadXcTTgHlL8p1FshmwrHC1EIou
nJwGf9gnwVfqxGhbcUgxLmeTJGPVvrHdgl7ayBNQBXSnzzfZoDa5hVVOlc8/BYzp
80LJfaAvXolKDgp/Y8mU9B2R1DHj/htuT1WN8gGZ/NFVnPxC2Yu6iusLZdECO34S
RvKCECKZ/ePvKEc1XaCbFKlqV5z+oa7AJL7PoBsWVGYTuTD2QLrE5bOf7Psf1Sqs
TxQjA8fYWXVpuQ+XvEn2JBWa1NIGm/gjBq+wn5zjHJO+ZnrzPgdPOVWIQU4kiG9T
qkoEyW0LKegx1PZWSYTvyyJEgTtPs9tYaiZimQ29F29FJCnenlZR8eglGwXy6RsJ
/s3kx8ApUGsVNP4a5GZLvjoD+4GpofdxRFqacRvWlM1DUwS/exIpHAaTUkouByjN
sztPshzNWMBy8JbudSZB8vMykA2zI+br0F5WuQptMLwk7BiQX7+oLGi7a3MOM9sP
TGGZ9y479mkruwRqxfH/P8e1vaDz5jUVsBAJyZMP0uvv+P0GUiJPVNeVI+oPGLnp
zwrz99v+uP2g0rmyQTEQjRn+J2D6DACg1Ix7AUd11iedCnuP6ZflJFkUvAI3enum
4gjgOwwj7OeWdYvhWG7v3gvHYPrFX0PUfTXo/5r2hzZlyQCDIAjVIzFM5c9u5sge
0cAKwuuQqgkfdUshCfEU8qVZksZ+JLYTCM7EroDLRS2djoLIKkJKabiiNo2KqIgB
t2A9BsiSZo/vwtxknFyrvjNT2W5A9NGFnFT0brPQQFvUldvytMmcwueQljQTrISe
D7tYznB+t4r9hpp2GUyFQ3brMtsuANG1qQC+Q1UQAeklt9Nol9fpD0zCBQCnjEed
6pIzajQlVmERs33xfcUYEuCcTfUZ09KPzrZmDw2rCC8zVwAG01sONrzAY1ixcrRW
ETf0c17nW7KOFNjQ6AqEtLMmEd/VXKvngG9hx3EMZv4QAQLQv+TLYpljKm3ZPeCy
hsRQQylFiA7pBbWXBgRNjv+sU2gxiivmN06xjq+uX1c3e6ADGHzT/RODw3QmODm/
uZNj9c4+KvcMNIQEGTXJ6IhleYOO1gwD4ACKp4Z9hnikt6h8Ux260OdaIaAw45Hx
iUeC2GN6IUpUQ/9pgdLpSjLizUMF1b+tpiFkziAvMwkjCvV4rx2CfioQVerlNkxw
t0g5uZuzF/nPT+2ryCHdsPKAfbCWphwSQTXLwu/Zm4oWLqSuKBd02sPh9kmXcobI
1D83ZrFLSD+0XyyPLHSk3Mat5dn6OL0+5/UA7CGLtku/bdeRROONR9BJE9byyZpf
QQPdEeJCOgrueG9kkcFSdbzTqGhSZ4Gf50p1mnQL5r0cO5WwM4N2qdXKne8cqSsc
3TMvnzudsm6bao3y4SOm2QKcUzk1ku9XC6QFhNDZcDBtV8qILTaRu510D450euiD
kb792/PdjtJmvjLPiQDmyhOK+BTmeWOMDzikzUEl8rSJZai4VfAkJHNZ0CKZ8VHc
raZMx9jMh4zpJA0xNqq7Vs120b6z6Oxw3oBLIg2VtqC+gyIpwQ4z329ew54ywDp2
jtevzaaHjNBkwiC9JADkOqr95N8oIKD+pWSmlOviq7TO5dnMlnIS3f5GLVasaIwO
20eseO8eoFL/C3/4emRtgodo5+IlhBwAahPK+N3Y94cdQUgawg4GXNwPhD+zTkGJ
+Hldrci+R7KR/b4M7ycbHufUW60n2MkRImZ6NFVm1w48OUpuEsg3cuG+X3JPLg3g
BlUzvNA2x2+pDl6ok+k+ETeRIcy0AWTIXRj1XOIrPYj05hXvE2IiwCATAYw5RIWn
a7mBNuaSIbvUbDaxIbWTlkya94dvrL3UhvDruQ9FaRHK1rJjxCocxIRFRzEKS1rK
QSscR2f25q9PnY1k0qY5Vn2/49l2E+h2vp6DnIRUkRLBzD+rCVsNMfSCTOqORP66
9kiOkS8M+f8JJOUZ8WGlAryBMpE9adGV8JPb/o/Wl+RJyl4CiGQVpxMdXnnj5x9J
4uGWfd9mi5LOdUxB7r2bXNrqzOwTEZ2wp1w8/DBxFf8YaCEBDMj65UBDR9STk4Ox
vbSwrDTOonv7qRqGtjmJKewNCmpskC8yStXYJVm4PMnGmtgBW+a4Hrne6g9U5Q67
BdcaQRA34NQ6Q6tCSv3S3rwtz1Eq815hdwayxPhL0hd5PBpVa/XsPMpycAZNMENN
bEOw2ZqG6cSmOWbDEUGSgHubwfxTZErfOfRa7VlG3uFOBNbtVXnrRXglsHQKWf5r
6nly/D3NjQ0Vfd8JmrjKuRdTtsOKEWTm8AkOVpOOzNP0AaeAHukHAQ4+9QXIraXM
Ig1HlMxjMWFGcnNdleiU299sJmsVUSfGoWsp50MRlT4XD528aacpm8YCbIDXMUcE
O4h31n5Hk442HsZGrMqRB7/v6y0e3/ywceV4rcWGgMVEoqWbXWjTXjvlLe3RR9AX
PhY1NHBKl0H682xTA3792rVvpimkUYpKWicOF9oOYyhw/r/oX7BI6QkEFun6quoF
c34DA2rJVJ0LsnFct2LqxM1lKpdjNmZHgvtjwH3JZfDjakgvCCLjCAcahOfP1was
Moq2nkER0kp4WAnuiPLkPWrSavKkCdt6A4xfqGd5y9blb5Ul/2+MRf1GLROteAaT
YvT+rYkK9a8rMriyb/pVNJA8zkWKdsV8mQwRNFCtBw14zOIROUYT66ODuFY3XMEs
kyFTO+Zk2M/95tf/9c0Qb+vLwNy3E0lFrgWqQb0n2Y3ae8l5Ai0Q5gk1KRQ7M+DS
SV8By/PLmeEun5acZqBnRAUWqig/sHjKdYt2pOrQ2z9gHe2S9ooeugnd529xIN0h
5YGPwlABY7p7ZE5xfn6S9ztdnFlrMLRHe8ls1+gkEu/FcJb/K5tZQKU6dGw9ny55
B0OZL3BVRTrArUcA3ZILAz7XTGMqkb05AkVvqj74hB8UboMQ6fdZ4duxxUM5HfA0
NF9E9tgL1pUNUSOfrZRnEDQjB1/XcmV2kK/U4QjbnjNYLOyqi97/EgX9JIaSbGUf
E1Cn3cokugw544oFD1hN0megDyk0t1vzgaLdG4danwK4XPNerw1OUujkkRbhbbca
itHcirsMDYHklf4FuH2FFgDnoY3T1pV0pOmdGs381fdy198Dp9ciEe34wpAOfvbD
m5V7sy34y2gOUFM14UrX0e/kqLHhFnYL3ky1dXtynMBHs5EmsD4Ztm+hDO9JWJ/J
NiebOtCNdy8hQLU/i/9jSsaA+RZxhMo7cDAb1nDSvsebpiRS4/e7WSVU+PvO3quN
PWkXX2r/3ChAoYccFj4S98dIxrUzU14S0pGJY7kNhfcMV9A2uGs/uIr6oLQmgWSQ
b+Y/yuM5AdAHpu57YiD/tCbRbPg6NwnKhEHGcZZeqdNa2XAV/xXYbwjshj3hphkY
3QBIFOqdiyJoORgXa1Sh0UPoh3QkcfFCfBC8wn0tG/L9xeIRmCkkfYv5UrRFvohr
Gj5xjMVOXFJtgOlEygoY7sz/I0BI0ha91iKYwERuUeWiTnNxN3u76VLJ563Fw2Io
EcH0DZfyun1GQiojXgtSheJSl5MD4bZI8UZVa7Jqj23/rE07E9NBFNnkA1bkjlmS
18/itSo+ZfILg7XRxRduPh5P5fOCm3ErOPKYPKnqk9qnlnQ5HAseZWcchYppTVM1
aep2/y1/8HCtgyBz9hMNXuUXIMese5YOp22heBf1gLkXYVHXhrYBhqGN5FMj8Wcr
q7LYS8mNn2md4VH5Zryc65Vnfi4zYNTNmYZ0wHejdtxDHfx0SEg+NT6BK0cEokU1
MK4vnJO6uIyRmJoPwu0On4S2dqDmzth94WUXEUBo5e/rVJCTdV2IH+6OLOwuN4dM
y+1QpbpPoROSHJ8lDpmiFE6xb9xQiTyNLqLp4s+Rle+GMgHJPs/6VD0sFGcxz6Gq
env01WfJzxShZLeUlh3C8TWEn2IVb4uCg+jfxpw41vj4PK+mvJh94QFdr3iPbvzY
VClBgdt9dr8aG5j8xRVDOLiNXUbqz9sOmHItmQfbVwtaqqmmyZjS4YVP79HeD8Zz
EjyGv9Oe+1SPpe3MST2zmeP/tqsv+ZKh0hQNK7vukvNrSCJtxLJeYUoszHCP/1WY
9Rrly/GBdRpb6IU4rFxNO3b52qn9UQfu3xhQuM25AtqDFPL0KbWMuE2+s9j/16zq
g8KXrEZm8efSdBSemGL4BmBPfMDdkiU1CnUuZv+lPV32bemyvzcOaLD097ceut/Z
PFA033Y9qu2YtjNs+jWfcPF7cdPLlgcIWUFq+oqP/t5fsbQ1VnuMh3EhJTtSko03
+RsghJ+XjTjVpcNJ/NZfF6W9jtxeB5jMdSBb7rYPwKKhl3HLXRlVCDzrTir/ln+B
1gb9NF6St6WErId25gww2ayUEB/mFt3rR2BdpWCjCyOT0JPi0guQ8OIkibOD2oY8
2rM8DLyWIb9PO2qMIFHxtlJQVgmmEzhfMvGWPx1SbrtE/+Nx7XlMex7XOX8yjXUd
lRLY83vLScVtb6UZIyCHwMePzOrWihzIMANidKqN7tk8d/NnpmRIUiTv+ZfduNQi
Qs2WFllLdJY9/aedHcA8QufSdX2QBlbcTca3vHQLBG7voVX9peoPWbBCqvCyjeo+
SWnIqaupU69SZeQTin07fNd/VBSQonqT7oVFgNeyOPDBnWPBXuxEBiogq8iaON28
rg8WWsB5Le18v80mnzMzf3Zs4aW6Ls/GBvI0kUFU5UCKeuQFGsUBZRiPPcYYig/L
IrhTyyH0wndleywy4UMFmDkwcivjpqpdGvRKqimmkC9DDvIKPObEG3M6rJMWnLpd
Wq3FrzheBa8Ct8KgZGJ2HR6AEc1X9NSGd4TlI2qkOB5KNxIT/n7USmIbLOR59QDz
pToa3OEIFs6hGVLbB9inN5owH15LDEVyU35UklBZgC9yh1fLzcKEUlBjh8oT8y4l
wwR/ZvKB3XkeqFiOd5j7ujAwOq865VEZogOXRiBSTfKkTh4xO3LJSPSwfaTddzb7
gXgCwMhPL91L18cQN9sdDsXZCsl8DuT0+9u04nuT/neSl/VJWABzjyw0JyL1pvRh
9llxaZ5JB4elpAqxI2x9AWPGKdGGX/lCWGQBtWh530Xw/Ef+cZax6M6ykLW0tRSg
Re/rWtIbupTmyZXAdgKC7tnXu0GPBi40dBMhN1ePcNOmNhKjfr1VYlvilp/+RiT/
QPasaLTkBhPOHsROWHpqhA2SPrhoy6LXua4ec7fUdN6tlzy0GUHzv6wEk/NAXO/M
xVmRIEXGAeBVaXORh99KHoNsg/bSDfxwt22kGBFJwht43n//+i9FFWRKLgYYzj8R
t2ZXmgqGsNR2SsuonG6Pebrm0M8XpJBrNVGfSLp3PcPyBttBPvYLu4SuctIts9bb
jcpodet8suV17yEo4YUq1CHeHDfeJVpjoLAmVc1VGYJNilu5mRRqLk/k0ikozs/6
6WnpkYzpSIgJfk674sVwdCg6g6KAd1komWnhfrsXIE2ngEFdwvuLESFWccukiYHG
ctnb+vBdeiPTcmvlOQKe1yq4LIhVfi2dCTUkhvWtZ/fJHy27yJDwKvZh+ySn0K5E
3UxYsSVMjGSP1oQjjLiKPxelV4I6cyIykLrRR7+iXqDhAeo2X0GGkmqaefIOclkT
EWEA5Y8CTx1KTWz0Hx5NvU/CRXK7alnqoHqM9FYEnSTFiqP2FrMK9DrPjVCHcJrX
xi4x67dzBizUrovqdktTzE2Nyc6KiC6a1LKq6Ikyj8peO15eNKg0R8FmYt3ojR8T
GqlOBE4cpnnEdCFBefP8Ytc4wUpVAsXpv9EFfldAA+1FpyEdOGfT4Zw7wyI3eVF6
JZyhoV5cUbiEB5SzLPFkXNUZ9niHWqRoSyT8kGyqhkAybUJxZYTmOwKGizTpFg2V
4ZWESiZRaLpD6qH1BVYckiN7CKtGGHXg4KvIbR5XIcz7psXO5jI5P6dW4xh5WK9h
TlSurUH+i5Fe5FPIGy8FZ+tYGOfFvd7on/atMR2JbSWNcs7CY6E8QHd3Q0ZiesSm
JFp7deMxlK/FI8pC496kqXm5o91BIFZfRhgK/Vf3U+LasE5qWmiOhuy/epdSGOD/
QbUZpJgN+56nK+MS42CK4OLWr7oH/aTFFVD43tLQzTY0hwfEh4lcGKT+hwvh06ig
bEPNbQouYbUhgAw2A837ygYAGMWD1Ma7qXXkPqQxtdSn7Q+77WXLMppUlRYQ7GQU
lDidxTeRrSJok7jL6MQk5PDvtmEWkuiozk7k4Cu8qj0PTAfyqtpzGr2lrxAqB6O3
84MKWjG4WNEr5B1qrpZujS9c9J7YH63VvvkBkcs+h97irUrnOgUd9fyj3ZcZ9ywd
ixKv0IceKT81ACYt8dq99FzL/VMddE32L6eOnOw3V0Z0/btsHh3GUcc1T3vyFIjj
cJ/2+EcIpmjhOjHEXd3Ol0io0MQzBxGLWUDeSJOS0oWYM8w6YIymFzG5o+nLY/Nz
KeL8ZgFzIc6m5cxvH84jqHTO7y/SNMt7YTl8k8xuWhZHFI/svBaJcus5Z6fXY4nh
T2Blnmpw4G9nJu4A5m0DALAsFXQ6l/qjOvkvQEui/JN6lFSGO8YkaflT6YXnA8Cy
iErji+Fv8hU/2AXFUq3fSiiRu7Y9x+YkjEQglBpfYjyNQJSb9xJpBaoWdcPXr6MR
vY9vdNAPaMPtDqks0qvnZW91ORg3URvJlOxcCjUqoKdsnT9sDi2/icfnJ3xOuffb
uh1pbNq56IJ5CdWajr9/h4RGke81KwwP0710xFKIsF+wr7d9Xgg7Y0mNkbcKBWx0
u/cWflo8FGfSKAXRlIckEGtOlOXC4G5SrLlAhu5WemO9s97nDDItiqIX2Gyaqnd0
A2zsYUt7UAuVaTWJsr6NvptpdR8D3akdJcDwY7sV0vJ2wjzjMgIDB4IlqdyJvEdo
w/CQF5azcImFTDy4VupkZ7Cg+8De/YJua5gKH2qxjh+VUmTvLb5kiIXztyQfbkgi
nBgefDkdQPF0rJV0WPwtO2xPh6xnZzWnoNq9iv3hcfwbDlRellNWLve7LAp2zLkg
rZUa/YtAFCJolNKQ3msTVJpjCfHP6nqs2IEBxFamnJo5J2hv1GnBueMB2TDTr8dq
3jCClvaQSWLlifUyV1cOCSbeXLWG/ZGKquza5z3FHisnNwQ/VzAuKgsnX+u14ROk
q8tB6L2mcoMsWLMOlUV2udntnn1qsKJklqKPZotSZjBTOOOXzbJBhSy7JPbKhjBy
egaKqIf/t7iGouJuWMuGiM3hSmEqrbBqrgw6CTUu1nzdMfLMGlynrGjFeEIxqHAP
RZYlZ/7F7vLNXTxadzh6rKUDkf2nJ6j37TSr7HNiURlvKaD1+XwzgYv+Qjtfms7c
Y8mQRGGPaYufQ0zskF2QgUTZ+ppu5xZ9/4xCTP/iTYvQF33XqF+1BkThfI7iAS60
rVQ2Y+J360DXjsiQoASNg/dinCxlMIDxUWvm65lLiJ/fYupXyYnxoDy587mBOSt6
r29N4HLMdGnpDP9+uwm2EhcTIMmpQ/oVNFJKHU4lfAPGwsmYxqVDTy/M0FUSPiNr
xBbTY/DmUMttyVjhGNI2QbuEfuNhZM+wu4HA4e3aOT6UfRjZ+5hP+7nYntiqJnw2
nZFzINqq3YmHFkgpNqMQYqX0ZVUt6gpRpXVMNlgr6yde06jJ3/C92jjN31a41KLw
bKa1pRguVqde0zms4FEUbdAnoSB3jt231ZirWihc0PU9l7QI0g1qo34wPGHMA2jP
xENImawMrzhvdVkTerntM/zDAEwW9/LDflDZRIJWoBxKqou/YCV0j/VqCjpJA5YX
v4+J7DKmAKhbAV/FJQCIrEh2sE6q68VQKKSPBFcjcUDiQMH+4MymbQFC9N9VASR4
wLd8TNq078kGoakhbvuC1x5h53ZY3/f6R4G61pH6SIrfd2Mx8mirOS4mgI+hc56Q
A1+H7LvDxukM/FAWSlKZysBiRfM/dfAcPZeQde7LtboQoYLOOfbXrN/IDlRtwbe0
OsG0iim3//8UetrsOv3ECXOFP46GPYsql6sPxMhHHeMj1kh+S9OnkwkmcxN2fSrA
pSs7apWHOuxB03PPDaxqzcCUwRH8wdOvFYt6np9j8+UP/POTW/022JAnPUKFzQ8y
iP9XruN0On5opzcOFfsUugKUOMOjyBYC7gvz5qiWn2mWAHRuTmkAd9K/RKZ8Stjv
dp6/2uOTlI+n3HZjdFltu8bd5APTW9wWc6SBKZhB5i12zAAh6p7nbZ2hJClGli9W
NfKjTQD7IrSJwRi79yHh9Am3WBWln4f6LjKMYcNarEaEWsScqElZPeD8bpckh4Jn
L2hslFkgILFtkmZNYxuVQ7xTa0LKaGSPnzkiGhuIvzGErxkHoj2gzk33AlwdCS1h
8Mz2msZiEgK6Fsemy7/lAYrtBdY/yuGxauzJZsudRzs6nDM2/nQQYMeVZgsxPapE
xNQ4WmXPYFCV/iMDjYkt4HfxvQrwT8MI8FpoXpUKos6NlEtF6g2ymRG6fpngrvQc
+CY5LM/1Qe1FPXUUYLHuvdeyqro8vIxeKSQHZaSaxUva0f9IOQqF6zqKQJfno+9e
TEr6HRpkxZQKvKlt0660hPod+/HzpSU6k16of5PEMoKYCdLdUbPPZffDQi0iQVYN
dS8cUP32iM00YjYYkn7Ww5iIHd/RlDzesn6hqlCu90CCR/XTKkM84wzOqGRLevx5
wHHHo3siq5pQQ8OjD1sCO3zfTlF6yATHDKCwdU8Wbf/Ckhxd0fo49QmlRyTEYu/R
ru4gp/oOAt+ERvIuFGSC+uXMzxkStdD48vlaNr+PIadaVPXtYXneVUqn110Kr39D
So/9XgwLhcEgwpLLHgmWvYpPFVpLZZZxHeSonm+VN/5zD3aAqJtu2X+iX5vIFSGs
FT9DqbMemCJVcktW09qMO6WECIIglswBc6MR3EQ0wtP6V/90ZnSuAfZVwpesC/S/
VTY2/UQKAteOf0XDPshRc+V98Si2r0ioy6OrPk7WLvCyCVHx3htrW8BLZYmqey2R
yEO2QZA7trZn4lCbhNDvUWF9Lm4fLMHOdiyK1eX29z+vZ/ngzdw8al63xxyB5JEN
void2nSEq3mpkdiqGhvp1dDAhezG2fDvXyExpQeNais1aG89kNc6WeG7cyWCePCF
hCMabao9IalHCze2ZsMPx/F8ve5oL+ihhTnsDZT32L/AgmHYVILMe2RujAH1FJhp
ch3xyJ7VhpFtNVU1Q/CQgmE56ap8QNyEVnPSEwyz4F7a9B9wLE0TnH7Rn4TnBtXG
6YBHdoo5tiWigUUYGvGm8V80baAijdpYtEeKNHPfm5YFGVb3mR2rMw2/7ebSVNqr
5g047As5RqlHWdKjd83dfGxxiFnJFSQ2IH6UnL7XNhaLBbJHS8nTwZc0YGDtf5tT
2gO4+sZzsjVjaCVCjCE831uYPl9Qnlr03B6swzFBvioB8msF539O2Xxc0092+f/G
+N6B1X7ohKSfd86cId3IK0P16XmoxrvO778jOk5Y1Ge4i0QW3TcOMUsxjxHGCyol
M/3DP9BGVhzT+0JijkA/M9GsbwBN0ZDul9IHno5HbxlcVGdfv0BXXGHRd1ogYWkG
bhyR2GN91ZPMO6K9XAEjuGB52nHueNiiXkuuaSxRoTjcniDxcOEWm/6dEnMGuhMH
+pMIx3H+LmiGRCfKxPqiktRAz7Tb1TT1ZX/r1O3RRM7op+GH59AJqBcI6sr+gLlb
fNUMDZFWXVpnRLM/dEvPRIyxVedKygj5C3N4wB0BQLw82zOgwe8Zv10sPKG8ivnG
WqBJ0wBy1G3g35s3/ogmHsL0MSogLLrTWquDd826V5pnNk69RUIPfygQn7tHV918
PBADU09nd3UNMW6K14PSScTy6/CLsoIapd+uheTjAlOqqW+yfGHyY1PTDKKRZ+d8
kZVb2zgi966wsz7IVxF+dYrOIM9lWOScbU0ee3j3sUQVDJEAaTDKYGpbzBT//hd6
uAvg0d7CKrR3I9xUcwHqTOExM8DcD57H/TpIfeYrS8wl4Vdvk8z78CdDxFFeG3WI
UvxIOoqduOt29uyodFZYftVclgyntHl8Prci1S8JUVB+q+HQkJXUCBH/fB1AeVl8
TlKkMdkNv3LUq5ZmejMQFiZ42I7YsijdzMVKawAkwoLauJjJwOn+A8UmnzlSTGDs
vr+nYjEpAq8O7n1xJ7c/CO1pzi+RJynCjGPT9Yr59Dm92bWdXaWAmts+gpmNIaVG
3dnxG/Wppxl+ViWpCDGQa/LNjVRMievMFpVBAbDVAmz+sKvFxvj3Rsw7ISy8Oh6r
qzrodiyzzrWhatuB72wHlMBvOoynLxmgDvkbzXEvpVDjRnpF0iZhBjw7p3RgUAXq
HOPnf0B1cfsM525W5jX9Yj8KyYvYu+bkLP4m7T/qoo/cRQhbGEP75t9rp/tcVWQN
g4WRTeizisbDf409viRwtwunsPUxHQ8XFft9VoGLW0fST4+3TxF78RWY+F8PKEnq
KUoTiHlcME0YWdaMmNxtfWqojd/1nO+Q10S47Rv54qeYGPef+quaQpCGAVZLrB+1
ONmyfHI80jM4F+qO/VrzQWHdrBfbP4XWG/rf6JwrNl2yKEIxsZyMA0naDnXyj6vj
9YMt9BQESfOdwUlo78mzl0MnjDLGVyLlbEyYgxGK3YRZ9cpo5FHZ4OaYs32pHYbV
Z9ptpCMzNHn62rkQO6GNeAtSotjCR20cY6wx4I0FQ0L7PwQIV40zjqjmktS4WWc5
DYgsBLfi2rPIZMmJkwL9m5gFgMbUYwhb7pihuu6zE9G6F3fjkmReY0NU81GAB269
h1F7KbWJl7OCRKLL20xcZRNDIo4KdlEo/yyDokpCPNZ3KveS3a0onwdMIVhti0yl
seOxgKEe9PV6xQPsKPQpzAlyfrnI+VJ8YIyR2H9ig6J8e0mE1jtaz5qGFWOdc4A+
uhEUOIg20s4Twa4cmtRQeRv1GLovRMqG2opN/27b1XdVUrHCSaBbP6mLyWuEw5LE
SdZG6lKNP6PJ49/Ow0SYKnXgChlNIBapGnVF1JsKDNg923jcwHwHM7rf91cvD22Q
L+RbIICArXBWzbax90n1nmcyCyocoCo8rqSsK72/ZsFzTi+tofnvZlFflQqGQnk/
K+TVheaxxPQKI1yLY0WRGTwirb7PO24JHTB2PuBWFxYG+ASgRVto+tpikxjbm9JK
7S5bBLZWCLiGkxNpCmU/sF1LHjpbGCHAPiBCEmHjUo2k/g4/30imRfhI7ErKe+eA
TYAf7P7oZ5ligx2bh8PLjjNRgT8R9q57rI/umCj6aK1g1MiaZEJOSaLMltix9Xsm
SQIp3w/N8IPOvmSCTGMXFfTBDcBne+HkUrXm9yk7LVypm/GvQ75QnKRNUS0EV0jT
+DRZlF17z4pdzFC4Fvgbk9ccp4r6Op0sMOlfKLVTa0SdDlAMkU3GGUtaMZ3qdjtR
mTitO1duI8N3r0f4BJuw5YqDtm4mf5R42MqNh3swcMQICJHmvqleDflQXIUWB+mI
1VOSzt/Yp17GzHMockC/XMasoLSiCn9MoKeNvNoQHsEv6UFveDTLKgDhiQO41FrP
cdMhS2eVog7tQLz4AH57SZVTuf/G/EMkSUOl3NqG4h86e5v8+I8OwTEmaOSlflGD
eOxWOwrTRba2/JSQe3L6AfOGS9xjhYVQ2dx1NIfgRXXcZMEzePYBwJSOUaJtYdeq
qRk5DZ7TzRsdWRgYystIzPm36dOCgEC4TJnzYVtJ1grYv0JUJye+54xH3Y3g/mKc
7xLQEDv64iaz2rtf6htmWd5eJbRVq6wtsNf6yYjdCql4MZBTOwcj6PDsWzCoB0Mh
RaZbnVJ5jGnA1Ikt2w7vyDGcPq2zmCrVkBjyFLAvnASrMeXzEQeNNvE/COGrOvbf
+V0voyfFTasDjgdW8aVy64PTknCVKuJb1s8H0orX7LRLGG2H0mKL6LWqaymAHcVf
E/wDcKkGbHtllAmvwReJWgOdGssuUZIRRLbNXKnvcALfK6BZoop3nhFlkmBYskE8
8ys00IZOotr2GMSf8ge9n7XVaG0CVzgg0nUlJ5SJfU884mUf+tRPYP0oMTkvsLUX
JT3Tg1gkKb9Sn8EgZGUkYHX3niOzKk6/TbcwCwSQ0XDDbIO/h/GbDxsh7KUWHcLQ
HqDHOHLdZ5jskOw0NGIWdjBU+ItbiQkrMTWvFRp1bbMhxjX8uFeUTVYqqNJNjgmf
1VKQ7UV5XU91obpGjryEXGGWBxnREB08nLyteCa57JBghjbItUx8CH9l8a4tlml6
nkxcqJ/bsLXooq0j7d64klIS8A9MturBdioV2XH5J5XFaWd4Vo/JM4TKVEqGh5OY
ixhcq8eBqPRy7vwKfX4chEn3brLz7A+EUImXtC/WGGz8qWIpAhN+juhEs/XH98jT
j9bb1xxH4S2eibu16wLVPypDXZ+ezclxvJtnUkZdUNyQ4CwNyovAH+9qMtTQBbMz
H75+lLWiJG7ASEBm4X0TAXQrgSxdgk8LWRKHtKCkp+27lDbwVQwRN1P2O8VTHZ2X
squ/vNilSbWFEsGH0OfO6PB75KFZrB0U8MD2u/r35j2vYS9VewI4fxvjHZDmOHuX
6WeKY6fhlXl6WsSOtguxIsnogH8OKle+YiTOmM26NaS4aGxat6Nq6GdGp+Q8Irhy
rVbc55yZGbez0+sbfInzpu/pyFgsk6d86E1/GlPLvPcbHjppgDZ+PLt9jZr4KiUg
Pr3RPoaZYzFqu+dNMyZMxNe+erM2Wibe9qiLhIphtdseCj3+KjswJ4cZojcm3OZC
dqKT0H7iUqwFaCa0oarnSZhyaX1a9b1iJ1BSKtFCNj3oQP4E4pw8f3Qql2pYoyV8
uZOeXhcCKMQYB/Ks0ybDDg6Z8k/rQGWNxZ7gJb1Bkgb3FZ/eYL+s7aEYCkd14qnP
5Bv4rEM3+159oThQXCM42EXZkcpNukzQx7DxpN63QqdveYPbsfd1yv45c4kTwa4N
4NqSyB1Uh373mr5FUkDq5bShiSwaiwsrwPnvQtLVLWQeGgEAPh5AtmWfentNzwe6
ZWi/2m9gjYt7+WqzAY9jcTKFxLjzgGTn9UazSdL/tIgqjSECs/OEBhiqhPXksOXp
G0LzNtHLoZKdlV0PbgTdRIJ36KophzzHJpUZsEK8097HyWv7XuEZ1UTFtc/bk9ds
Q0mecDDswR6UqzoAdf0MxlYzXgsP0/9IKpjR+WuYbqAjSIC+pe039DWKBm/fhKPD
lwow5tFu8IDSBBJZX3g+iq7GUlY0MBUasW3JCKF+UNQXal2z4CMdFI457cHk7WCe
ZmZmEf+rHPWZ2SGTlkFPdFtrB4DseTyH/5oqJ/wFBiqW7+IxISFe80HiKlHSbZIi
UQF5Te9Olpo0Te7Z7HhTMcrrZAgCaDBnCoH91RBM4njaY9/d1lwhXB54yHfmQSQi
gpRX4qc8dgLo9sarcvu31c+dEy4ICiiCHRaTTOBF1vNOcW22x7Wq6lYR1FYJmRsf
ae728eO7n5IG4kEJHsz4mxaLO5Sqrh5grCNWpJteKHWGTKJYFlPHBmtGVI4cLAiB
5bauYr3kK3WWZ70FsEXZqlsDST67JekNmcGOfMDaLfzOq/RW3WuwpWw4Xsz4hwCz
pqTex4kysr6RrrDHK/X285T4K7wCiFUVbL2ZF2xJzFJSmAkCsE/hXtZaXIEtWJx1
G/je6rqP+OMeGcplaAV+YS+A+H2oWgtfyz6hIPHl3ysTmWjSTmklCErw83XB8nwp
/P3GVVYWKP6cg5OyfJ3M8f0lRhIDJrnp0lWfJXrDOimYmVl6bwOZoNp8hlXlc9Vc
+qKxm2MLI3MfhuQdHIBtUadLCL/EMxvVLud3qyA7I1VGre7XnnheUz1GR7op0fO0
BQ1cYZ/nUKN6EbEooHQXox0Y0jykm0aasqTFG5/waFRefFR9+hlfF85+0p9GXFHf
iSFCiMvl7nFvCsfPh+EJzWG9sQItCYdMn2/wUiRO+4W/pZ/zI1HgWXxcwPjbBhgt
yySRDef1M7KSFr5Iz/wn1gMlyO5oU9QfJp2L0/XmA/65XUCIYramNy1OtwcQQjZj
eY7MgRhMbK4GW3z3W4jZBuxh+zsvjxbPfaOUTl3gOirfNbF4lRjm4vjXNTNkfeCk
8c8Ro9BVlP2yVMxwBQ8A9XB3MN4biGH1FvPpQg1uiLZMNFNc/jsklOoHEDKY5dpD
4+lfat9+2tt96nYLuk3uFgvW7uMs5Yvtk/HKc27oYnrYcKsnDyHXjj45Oobk6Yxr
PCnjA4I0GJDV4MKysKAFerV2gS4yqTQtBo+Nn7wwHklkA+bGN2d7hBrPOTatq0X6
mzzzttqk7udrFcG2CpcVb8Cth7O7nBIdi1Vq5fuLhyMu3UbWnBwtw49+TWUNCBXO
YjE+dRiIKRvQEnr38sD2Sdrez6+sOl2C47Nzc4R8eQJnC6PcOE60gZpewofxmZRJ
msXJRSacopJ3h7bdIFEW0VRkeg/Im2+UBLObFVrjh1Uaq+atilrM/U+N6VLVSA/I
gTJMkn2U7W+gU3clPAzR2GceQC73RYP7L8eListebj3KUeTsk3fJ40yiW6haYnyT
tISlK8++lC5vyKD8KwEE+LE5W6xsL2UGsrmfCGNFt8OxxgYjkqmM57PcgQVQYKFY
VVguRFpPIgVC2wRa/Fxf/kvMDcs+Zv1oQlmWpAJEfS3feFurD/gxmyVSgrHSecDj
kydIGdQl9/NGEu7YpyqJ5OkDG2rGNLylioqjePE7m6uX7t9VjAHeGofGfYCDxsuH
kOvP+IVbQJfaQ34ajQTselKZpNzdaDZVn66GcgXJT94MuPAnD6o2LRAhrECaBP3a
q1AN3daZOqzSaC3TkkYy0vWxxMeSd7L3jULD2I5clU0ytiJLUxZBQoTzqlrT+I5q
xSAAL/qzoLv0KipICeA0DLrFAexuBospnt+HBEoSE2TjyRzRK71BsQd1abQ8Z9+2
tphnS57tS44BrMzxNiLAJI0Cz2EpHog8XNBAdJRmSj10hqmufL4X5JVdEmb3wPGI
POveWpYwHjPR65Ckd74kWU7mj/Soz6SAVltgjIeRKZKr0n4BNeaGKzSk28rXairO
MR4IfBnM8RGbzWFaFRZH9eNtSPvyFAQ+zTS813Cns/QGaqFNsGQO9gp0CjpjvfX9
/3pIo8jpUBUDtnhFH2vlMWvZ8yR8E4/npmQLF6576BwZrCZi7dbHNEX5tqLthvvy
syY3KIpjR0tvp1lH5hlv9kjobQnoydeXBYhxkGoe5OfkN6ily7ciQ7JOAw9Z2c4J
TQboZZOS6guYwVAVn0tboKLsbBl4+edRQS4DETyKE6mc/psnavsUGWbuE2mTA5vI
dgNfJ3Mk9Eo0kl5ADNbwopR0B6vClM/TcMFkRd2Z0DKQ3duy4PphY29fZNgg4vug
OKrhNsDs3cyNcYCKYnshSfZ2XyNhI76QHYEmubew4QYizQyNO/Bf8QD8g9Fa4grn
ZAXngcmRCxIh9IRYAHOG9z91X93cZ3/VNJI9tpFWEXfVwVvd/dA8apOL1IckbZJQ
SAIxf0eDEJtf4LRxnCmxnNGSa0X0pRwBOZfDQKidv1HuT3Hy78cSrAWD49dYMWUd
D6nH6LDlaywi/tswx4Joyj8xRhm+F98cMIGJveUZjt3s+qEeKQ4ZodfeqrX7gKI7
RlZezlIdqDPMzOigu2VKP23sQEz3suil0cZYu/dRwr3ptzD1HZauddwSuWJWwdez
K8elZmjiMKzaDvd/ePBSLm41yYppr4aX7UgjA3zasqFM2s49wWtwGXmfNgk0ljM/
jW3J9bCP1qI/eotnLwkkl99J2JOQmsis6yTFA6IvLeFaFnAg3tHJqHfBhsi4heF9
ts/BZYhryJFs1Jiy/btAt/2IpOmGlnGrcaKQgykoreO/ndgV4yQwmexlu/+cx2DU
H1Anj4b/PbriPcd0/lw7qkKYHSZi6v1eN1F0UkUrNquw+yhwCJZFzDLfHiuYBRWJ
A4PcWp0RX8cJCmTIIEhL+kjektEcP9NPMA5hNEHPKJltEDdbLVXiFQQoXJS2opnw
eEqp4Otabb4y7oBrQznTtqCmc9PeA4vChJ3CWxL4TjTtOuWRXl0qwnkQeiKIRCcq
rxh/HMgsLSQY6qBQl7++Xj6coYycVsJnrcEGYHpAcfaLWoV7wzkuW0n5cZMc/ZK5
n+U2q6S4yN6T+mTRbEey6S+gkl5UBgLbmG5ito3GbpmTth4LeSt/C+tHFJ6BMmAH
1uZGIA3NR0dsL3Uog2mMUpv32kg5m0jNX7Ue6YYm2DBI8+Ic4+TUMbDJjnqpYbMw
MbVmfieE73/AIUSqQ63+7XzOTUHLdVdMVlkyXFnwGDRaeIUJ29hARduFNFBjl7NY
Ur2/sOtQ467m4j15kTSREXC8AXny3OMNxs0IATo6dEWC+BPXbDnL+8dc84cd5Arr
aKGfXFbsVi69bBHl/5XhcToq6JSpKmYb5amVAmgemDeCv3GmiEt36IW3eu1xL5ky
8Wjchb4yB+O5CD+yCzPVLfxRYi69oThh2PzhN4u8GqJG0SmH2jfdYNMQc6MEBX6D
Db222kGoqZItBlUn/zuxVt/igwL7ETpKUTUKpUD62q2GUKwbWRTR4klOBLjQuzxG
hG5h7OBUUhquy1Z4m+sSORAJjkW5xvn5yMtK7W5K1S4uUUsSvNR70KOL3r8B/lxQ
zieuIphM2ZJh/YDyIFq4Q//efnUHNjoTx3k8Q3A230We88gyyiLPhry/jIhRL1ps
ItCplZF358QG4tzvtb1PI2zFmHgUUQdy1WWn4gSqQSd1AXPif4fQY9Fmbk7gazrz
DMA2bHLGRT5AR8o+m4smtFfvo+aFSIWNw62VhLr3kpecXZEJ1yT5W9C7HiGT/Mys
2hfsV9FzWLiD8/7HVhHnPTc0/jLZsGmKaU8tj2CREZ2plpNGHfOIc+LwEUfoZacl
/lZ07zz7xyBUKxcJGcxnuASCLCfYcJMOOC5GOq0JN5OrC8+AK8EbKKnCGst2i2zK
nld6/c5P38rhajh0eimWZN1IO2XN319k+AQVNmQX4tTkiP1IKa/tljR9utAz8dmD
eSc9ILpI1IlWFm0ojoCO4mohohMZQkf6/zaiChW2ukZV2lP+dbulgp2xbuyMEZqq
H5r6Kw0fPhZPGKj2oYUWVqIrABEn+fcmYyTsy1t8Sjw4qrjxhCPREFIm7xWHMDjF
MxzsGr27BNhovdkh5zyWYqHPjEfC+pLOTbvl+6mYdzvqjGYa6WCoufWBcNCepGKQ
JoI8Qp4lWaMnsBvno6ZhpDpq9yhCem1KZ4/ewmXWJwxp1CtYl3cbCsCWgXmzqPs3
KaZXbuAJTFUuyCotlVq0n7/XC6OmIZwk33TNk9bjmScyJgN7YYX6Borl9mZU65Sz
mVNeGf5QGssezOfOzGho+NuSMwDt1e7u2LFxScbDsBJilkTFoWFOkE8bFaikkTMy
k2Fud9Vi7XzGfLxGEro6a42r6xI7hhdxuo5TdQN9qIxF3lsfEl+tETeCLfFR4mYv
vFKXpQXnXAFSBQy4piyyzWexuvaKG+YGxEvb3MPnlOv+TQJZuW29kEewaQMg9god
z+kWXT6qzmdQLeHh7cZQl0qjL1BcGhSH7DrzrZO88XLjlvh4afyUsmXN+jbnoQDL
HnBIoP8fuBxi6xo91jPJVL2z1q8tpwJ8IRx8x1Nh5dlpBuTk8qKM/mxRk1+j7+Jy
+bTYU8cZcrm7lFv1EGqRTscnfPcC59954zhgtvkOsMR7WM58iuGg0k4nadU7sScX
Y19q61Hui2865zUEm/wSmX2yBzIx9Muipg0AF/Y2RpSgd6oXo0YiL89smale4sqJ
zbI1bMy0pkcNino5R7nAQ69SF/LSJ1haBOxez551xKuSowhwcnuFuSm7CrjnJhg5
sVxjsba4gL5wY8b177HCgbhihvBE+rJT33rdYpSATpALng7pbu3v9Sg04d3ZODDi
XGGYmLCCQkek4VS7RljPUhYszIaty8GVtiHN7LInHOY/yuo+oNNUlUb+HEDaT8nO
i8U7dwpgcqf/5UfWYL6IXvqEb41Zht8JylVGIkankSKlHNLT1MMDDP+zXIxnWS0P
wsjeh3iN5ZpImyhOyzM/j3KIvPuVuN3f/G2h7E1fBZkuL5IsuaEgzLm0ezkRm5NE
nLfW0px4NGs+fhadengd/EF5+asNreTQDE0IzZeJ/doIFMtP7Fi7XnHEUgSDh30s
Oue+3j0py1MnK6eLgAMUoeIL2D7cv886IQDdD9aMG0zNAPtWUOkmbuT5TbOmcGtv
WE5VVLxNo23zaYaPXatLIE9lF6DP8GKxntxC1hkA2e4MGMhyj1qW5//swxzIEKAr
NbzM6ag/98h7wrStQ5k1LzDOPtM+muPcRRSwt/JeE1vab32sID06r969yytgtiyD
R/2a+nxVOSgg9M2Lj8rrxZZvgzA4t0CXnRVzKtFVW42b+KpE0c0im9FASt8K++jB
Y8OaOaz3LyYpVhXv9eePKT7ahT6vACaXMvJ5gnMtsIh6NXWHAoXxg8hciPUrWtkv
AAO+Ql8AddYnc3fvjDuhzYx99ricjQeFp17vAl6yZTpR+ePYyfuYtC4MSkCu5igc
ApRrQaKO/v8Yi0oP5b4ozss3TVpPF/vGTk5mnBi1MtCe+zf9oOr8O5Iq7i/zzqsp
6hWpuMQm19h7+6JESbigmGC78WlrDXYocOkOwEt+wDHRwQgFHxXGULVfSJRa6L+V
HrlWYhz9GVgGmWfXrqQUzRLItEtaJV9LU9w1Akbd2be57b9XHc+vdsdI0JJvF1Kj
0WZQn7MQl4JK7MeXNEVvaxwMNSigelhin79jpxTHbfrCQzmNVm4RQCr/m8a8q3GM
rLLZ8rpy36FOUQRdSpevWRXWFsYrF/K+Gy9dpeIxTqpW0NJS8wqBLflVv4ynz7mM
sBAgVv433n23Zv/dcGGxoj7TCyCCwjV66r/LmJZKtMJWTDJK2ikcDgEIHlfk9lEU
tnvKLdPEI8+xrSPa0xxAeMoFyRrmYKbGfibZVnXgshCteVKz0iwslVWEhZE0g3E9
DRgCbAuqnW8wsWZqVRgZtUIuAwtE/2u9uzWYYOGnkGTyOBIvboVOLGN4SUQyoayl
/PSIWMXv67HuX+vNg3pkK+viJQW6zAOOReez37VAf4PpfSXMU3KFSQDtYofW9KgR
5kGVxTGBzdSIIJ0+CIvE/NFODrRiFxPJoRIvGahFciEorOSyLRe/PbnUTRziOZRi
EC9XAHO3SuD3hTUE8WeB4LKr4MBtz3oposF08S3Qxi+7hwjI0RgaIDcM9W9avvD7
t5ZpUs8JIsDL79HX+x9QAbk/yFQKoQI2Whju9tray7sXC1Wux9x0BJEeQsJs1+fB
whRXAFBFKtghGoCb5S7os5voiaAnJf8EWCnmiNuWa2QomMSiyVaR+5PPeLIpir4D
l1JDqvzNnf5tgXcSry5JDKBq/VwKSqRFIY8dZJ6D36nQHor/LhZzWli/xHj3DPam
ASvB91YkYDwlQbPrK2sVa2mEHAtKTuSwKzMm3t3By/XD5I9rke30L2tGtetkUFkx
DDD2DOQC/vjiXMn0JlHsUHIrBqgbjx6ynA2ODmevkZdUBgC80kYIkRXfZYWTxAXQ
PUrJS66Ct8XPM5suSm/T+hOAbIRzbkpFiip8mkgVNnGWOBEFN4COccrb+Ccw/4Dn
6daz84VDNJ14PChG2dyWROS+FIrdjiBFOhd6B0Lcpa0TF5zegD67Qbr9RxJjozy+
ZKXud/W6c59GUQ5Yo19+/w/fw/vssimwafbrqynGgF2ZXSGFH4vooUvHYgV2PF1J
CRVX81YqPmxYDtvoVv44nXI57ZfIKScVb0XYapiLNUpO3qn12/HgAr6C/eAMmzia
8BGVqeWk6XrfLS53PKF8uoU+Au6tAGS87LfNcclGAQm6ygQgwk8lIl7y9IB7J5BU
bAhRP6fKEY7pWWNgWHzsXuQsrxCdr+00tmZPmZMq1PzGV0vCEp2t/8WzM75RhLP4
qve1ZZwhdurhLHfirxz102C8Xv7XKcjUFJTjAAWuMIFWOe8O/6ZtpYCwyHQ5Ujea
uInSNI/jJPLxVAf2SZM0Cpmq5mzzW4mNRwzBcbHH6kwnx+4zOqbR+v17qJGcVaL4
YN99MtpO+o0V8gwZ/S6k6vRmjpqBIrle3Alqaacbp3QHuK0pouGJoSKJXquxEYEv
0k5sPRq2x+QdjyTAqsgsaqOy67cmNGuLGnxPsBdecC/fm3NenY+9v0B8GobZhb7m
nZEqIWgEJQMFd5AZhZ16ehkp221KExYC6x4ucyeD1B1n0ZA+xcCi5i8wE6etT3xK
UpX+CFoYThAxdziSIp0FN863WRviouZ+OW6+Ls7TRGxk6IA/cuOyUi5Pm7PjRDEX
J4IBZW9o/+8Dqp1igpB2SzbaaeMWyaeMDpXnEZwcuHotBIXl6Ae/qfazDm17tF5j
ccdxq0cYNZj74+tKFcnNLil0fri2/O1C30DvtpohuLExEX8eAl1dx3urHDEWEnY3
f/QZjUIN5EaSl9E+iv0yLtIHZXd8aZw+g9nHJvfXBzwhbvUpJrwO3BZEjy4wujxR
PoeiBS+WVwd6w2OXQmlAOxm8zNHCiqyhcBx+tiEfy8KkFZ9/WTAAUAt2esATAWDb
I2f2RC+7Frirywy1WtkjPolY9vU3n67CtngS0vy2xDp5dCd1Z7XpGz4kGItBpilo
M+2c1bDMW8NGf33h3BDRTvUfhTW3LF0DpWfr3MInA5UoX/aLIB/2Y2Pns2rUcd3+
rGXRtkA8vEfUb4/RAXNh5VdTlifLIn7HuHmdSTcr5KYx18N1hnX1iFzd9TZlCguM
2upVd2BwBFl8+ChS5GUANyl8u/vO26preWYoE9nyYkiczhL1LPEs5EEDsfx1ApXM
RDC8ffR48J25vTXT194dyNsCDwIOFStHV27H51zCbw9ZOqjAmIzFTrRsRH1iWiQ6
hpwnDP1Qbdw7nNvy0MTpJHK9+yFKLzhX0aqPEUvL86DiZldkqp2h7CLbAigP49IB
9l/RbjO5bz+WO9eGZzC67DuzaB2olHN4zatn4s01oWZ8wTzNnIuhgOPuCQMjvM01
4i4P2RMp3du4rokj0QMaD1CYWrIzgWZV/s26Vs+cWqhhV07NZQpdJ1iRH1dO5Kvc
s2QYrdOk3wKdf2iw1LKOQyndL7LSz/3jXm4AF08ug7Ftjlu8DZt7P/PwJj4+QOh7
pCTi8NwqUvcdliZ+fRQQ3v4t5NDYvM1pjaRauqSRUslC3jhwziGWJF34co3NIKXT
NjyV7SB0mM50+UJ2nKm+Nv3gx9tEuVVo5uqGJGsRCMxV4ktDV7L04FdZaOYzDWqi
7Z+PqPCDMbpuH/Bw2ju9cLwEq8p3nxuqJmWB6gJFL7FR2Q5fO5T5X7peKfZtWfzE
HsDU+o0irQ4PBmf5TXW7MT7FrAoQPIpZGR+cdXdCcNzmBizj9rXqpVHibQht537N
J3TCkPOHMBoPQx3wKCxVbL0cXxhO+ceAQghPUX6LDjkhAmibTHeR6Jw9d0xua05A
89IiUFj2xwAssoHCyD4PG9EnqAwhg01lI/2UDttAIxJDppyoi2ipuAYQvXvMRn/s
42HrMjBrrAXegdyDY+BsFLC6tEJCGv8pJnWYUpcrCtQzOjFYGKz47mzZBgWF9CMD
Isixiz7B3JdZBCpo33zxa/Q5a6tRCznIbCwLsFh/KQFCx7B+/U7JRmSYEtlX7G3T
gR4qx2y+2rhXnkfKFD5M9+MWU/JozcdKjdeaqGBZZLo4YlfoMcjsuRGf4iPchA01
kcv1RE8Ezm0FJH1DBKCwzGnP0jG8S7TS0KPpdaDBDsRHF21uqHKcFEFe2evupdFS
0crVMO+MiI/foAwnzeO5of8wcTmBXruLrzzWn57ogYViSZHt/Sfoxr/R4h2gflds
MU3WLAcY/dyK0Uu7YtKg7z+WqJq4MkE3zsXM30sfoZyZiWPPjqVgmR0ox2L2ka3Y
EVRJ8ZUMsqmsa4YKCx/8NNUuuYDOPFDaRMMbb2f3ZEXYzeiqxmuFStY7Lix9Q59R
Aj6O6cMYOdYBUatdbidlwGCuScVOSkQ+IjuxNT5vU4Eqms0OnrYyr2aSnt9scmcc
LMZzdSdDx8T/W0/BlR3sptqNcPBkc3p8vLSLUafPGazNFmsD5iLhVsxfm0qMbCDP
3HKsSnrzFrUFJd4z+rdO3q1oOA/7n3+kmvocgRl4wRJFQXVZ4e6wyqJE1sT95Vzu
UFjdXcBs2YZkWhPScBLdEXVwGQt4ruRFtduuYyYl6EcO0V1M6pPlcM1zFvUCWzUA
FLiGwB8IqFVw+1aLaz386dxtH0i//ejR497dgv4MzuxVdSSM61ljnjiyHdId+Cwh
KpzlY8VjIYeu/amVTtx4am+XJb/78zlnV8Gu1MQEmCFf3TmTjRrmcaTojixNVzow
/OjPHiJhgnd7S3tWtvsNlMo7Plx3Wk8DbLfkAk2xlB5albq+Tmgnlg5q7Nxi40v0
EEJwXkUQdlNa9wMIQYhNl9pBLdlgTX7I3xWHbsqk8S+wBfJPeTMAEPgY0smj8DSD
XgsNyZsFe5/0YOBZnVvGnZ6WnIQl8M7N4PYiLFPRnHBbE0j74K/n275h0swTA4Zf
zgOrknFdOjz4RQqw03VAKwOIjj7BVezGkJ4SoEkOPQvMkLPqWHmj5cRcjO5JSaWu
p0rIZw3YjfYqWlm/9gqhrXvzf78LCtmcXScChIrIsy8wMv20d0+RwDhMFZ+B9ViB
aaS0+loTUkv7JktmNHQsGUwsxOThbR+d/sC4/O9kJosJB5TVsJAwTmZZ2oOq8FBB
euQ8e4lJ8Y5daojNrr3NHKKW3zifV8bAj1EA3Cw044vhvlRzxfR2aNSZ7Sm9fPF2
3a4nh3pqZ1kcWenT39sytaHQOEmdrC7+VFyXViY6ooreXd7No2tJgOuyg4F0Quf1
4eMDd12MqhjCuTX2ZseKjDKN2XEgfeTEZJwchs4QQbkyuIeZ1WzygkPnXY1UJ+eL
xvdOaObQuJLqMFi0AwIx+5tuLl2uqTACrP3C91zgg9CsooQnRb4LpldtKXcaEMgv
F0UqpTZh9OLEV/FSjVRgDyKf+SKMCzMAPMbzkvDGyya4w/9N8tEzUSUlxast1byT
XZh2N56DDBGTafgARAg6ex5UXF1i+7xRZHC9485gsDHCP9PuoZA8VyPIEAZXcOiN
1ojBc/Q+JI1HroRcNdOENTqf9jxZP68hvlnebV2/v9F5x2AzhSw8kJGuRTBQDZEn
SnsvbEDpa2qTT8BLETIweQ+vXvEq2X5NBbSROEwscyyS49uU3C6zAfnikGnytYyk
WUcgJPGBu/qNoTmkS7wgwjTEq/EJ5sF4KFcDAz34T7IRirbNj+sGjJMmoBJfj+J5
bop+SZwNfyACmc+ijz69AaUM+5b0JngmYH8fjVxrCQ3oP55P/S+CQKJgaN0Yl0xP
ugcrDKvEACJN9DkXw94vryDeozbb1Hhr0OW0XGkHoeCcn+CdlyxohF7TtpDOSrr0
YEOrF0xndaj/62dFfaV1tfSThkXm6G7FpXU6XrvuEMM7kwf+HmSAWPe13I7ZztL4
DOmY9DQHun3TQjv/poImzGpsy90+4upIoenc2Ytk+DikQpjf2RWATS0sKSxYSolA
xCHmGmuVY+TEz6LHO5Qu4rjfq97M/dv2guvWHshY1oxFW2+8Z+lqoNkc8YgdFoex
dq9a7CZVVrwtY84DqDoVymuueodm+Wv5o1bHuwEh4I/kCb7xwEqW0Y/gfwyM9flI
Oqz9pdNX0Nt49phHb3r5eHUJOSxBlgYdXsWP4aulpnn7+hbNcxPw3BypeQTLXpOW
NjE/i7JDrdzcYkvsdAYDVCJFJtkltYWx0ZMsB9sJjdD2g3Txgw/VfMst3buZir+b
raQ6z9GZ1CLTRgxkcyqQfloD+u9EAt5ux9WzYYnUpLgRDWXeFU5TX8312W8LP7Nr
lYw0k0GLgARQn+xOd8W7CWB/BtuA3zeRimbHf5QIdYmlsaTlWcuBmjl8xRETQW1N
2sG3PktwSclLlGc/CWB9q5dEX79Z+iEAf/tDoyYi0zoX2cdDSP4Sft0ILOKsXuM8
dT2lAAjdR7xegzLj+odnf0L1Ita2DNtGqCJo4WKlC2is7GVJionMigia/FrndPT7
iVWJgbiXHG6pYKc1lK7o7pSwATUm/hLBmKia+0uspwEnopw+TvEspFriEXCCHODm
jfgQB8UFRAIIuAHlVs6EDioZYye34BGZ1xQgcfPX88fL+SSLG6KYLcu2RUoy92iw
nkJ4EUh6ayz4DblrGzjy6ZdKOQEFNGTmG71+p7pEQ8zr2WIThi2LXRPSWygAUBdx
EEi0TzLvG1cABUPjKtctRI4N+fVYKLx884J9lzPeNH3z0C/BJF6GAHOBRoAhJ8N8
g7jbuLF2CHxiYbq1IEeQoZwiHYk7C9h7hEWKFyXX8xFe6YYEwEPO8bV8Ch71QZ0c
ECFjFaSJkFPrJIQM5K0OqdJ9MkcV8g+AYgwDPGLb26H1RUjjg7t5bGI/dfEIV2Eo
6FKHo+DWw1+bajq5o0EIbfXr6DSczG5mu48zmq9G4n73y890BzZL6k82uCNCeg1V
ejy6uSF+Ul3y/rMad2nEh0ApAwqZNv4Kpt5lNGxKIp6wG8vy6VE0WBHCUyzZHX+Y
tEb0SLVZfhzTTs2O0lqZ2pOAdzHGZ0WPxgBb7+nMyCeWj+AsLk8j2fWSc5MlwsjM
7Xp2amoI1dSJX8ev84qHMG/JyPoX1JDcI6X66J2IuEZgS+cvSKvNLQ6VvWxXyJLY
uDyATlJNPds85oQ1NJ3MjedQs9Y66oNOKPAv9Ebiaot8Ig965J3qg/7StoxwP27v
epz3IizPsjtetV6uxIXtM3GvJ59L7YAYUvs0k0Fdh4sUjf579TauGA1vxm6t+/tX
anguwrqM+Mzmtm0ajbz/S5sav76YcwU6Wqv3YZDLfGQ/8Vgu1yYSGtwBewgToUTP
491uLDk0sp48biy7T0N6qD/EDHOMM9uX5bfJyqfi1Rsiayvl/8CPKa/+BaQvPhFv
3odMkyg06nuu52SXoU9cbyU8V7xWA9Z64ac0Kq9OclTvv8Wld912qXiy+zBKjNvQ
25RQ5MmBtskHCG0KwJXHjXwWosA+zN45UmJjJmth9XEP4FJTBUV/rhSgPvgo8AD5
SQkwDsQ/2I7OSk7uCL1zPG/ZB01899UrTmMf/Vuobi9FHesUalmyp5wIqbB+OUCG
dzNUL8lr91LHU0MYei6qttLGrRZHJoNoVp0stNga8Liaf9qBbPefDA0p3FjwNJoD
O8oBFr3WXEKwBTs6NB+1Fx35GxcX6acZr3S2aktAduwJ5rwL8f1Ohdjo9PQ/HJkK
hew1BPVwzNM0fKIK0TD0hM4gP0IfsI2PGOn/tShNOSP9a048PRUMvK48eeSEc/0I
2+1y1LqzK/K99unIxy4Obr1sGYtoAia/s9yGZEDi192xTSRutQpxAc+aGZfrjHwl
v03YsBJhqzcyI95QoQQUgH/bEJHIFMuepq0g92wkToo2dEd4Wz1lflFyble38n6N
rFd33xY//pwiwqAeySdo+Mq3OQUPzEHDREg/bldoKxQzzuZ26CZS0LJgJZuQU1VM
YO+0HuVPx24hQo+MR+2rgPQwpzMPc0c/ndJ4R+nLg0N3zVtNebcTO8oXTJhkaxRl
k9YzY0CHfIEjkdYqBEVk4hRXWAmWzu9oBtoqaAjzzlgjT1d0USbySwWOGsJYGusN
FveQyT1Tg8EWza3zmI32uWzuzbR5LKwFymtA8Wi6N1a8gUxDwQBK8KkYp941KwPV
NNcjmhHxpTwDlnjDH1n/vA1D1sr7udLieOP/HmqMzQUmhSs4fgtILtYO1zdn6PVh
F1kFBOu9pepE111x6Ym3vl7ak1ChFy+ZiMKibtPGLjX6/mJtpZzv5krEjrAPRIg7
gI9vKKEUeoarVuLdwZwJXAhC6flqt5/hxJWDe5Rkl9cWarzoyYZjSihWnTQ3r1km
Rxj9v6//6xKowE5B83ooDsjhOd82etrTsKfBCPKTz6r5MiJdzGjXvC2JRmp7yhql
/zOqnaCglv+MooRii7FEVsw1GtkyXwYZlPUWhcDN6eQ2aFe06kJBtZ9rqURNHh7q
FFrAm41jPh2I9JjkGKrfVfdKDPTUin/E8gWqJ6B68HWwzCC6nPdG+sizMYe9rSO0
haq2DVY2GE5NwbMDlV6ziZL9TXU8LAtGKQWbYkCy68xo3fc/K9GRrJMZgxOAgcPF
+NMbYY/PzdNci6uDE/mR9uojaYb0MeFb1MI8CKwZCNENlALdwWlJIS8W8LmJEo18
YpRH/PV9dEiMPf8yBGffC+ATbwytumY16BAiDuoH+qW7Ywc2KCavT7pUCHQ1KWC0
P57ngl5LqEX02wNREKqabDX+Snrg1zCd/KJEQPfPi+Pma5m4lwuh91cS3eO3XYlU
xqD80KJgxHZes4Nqp2P7ZQ40MBUcUp2jsBgDarbc7H2u5wbi1Id5PfBuMuRiqQeA
hpnlHRyH/h7xUrNP5v0HHImfMBgaqoV0bWJl6tHpgAAY9CgEJ47LG0lv6Thvcjyx
75RdPX6jGbNBfcx01WM/Efi0qLaV2P+IV/2uW4lTofzBjTPpWR+2JcEJmaJDxZCk
TJWWBKv8hG9OvDGTXHw7AZ3ItkOoPHH65QylM+WdD/QcEdP+mWcFtf7apzo/IpG4
qCiHx+4N4Se6bV2D6GhSrYcs37AjxAnP0F4xO+x7O4M9BstnP46LX6T5hwyLhc9/
SVQj3k+MVLY2T+EgZ60+D9GWkOyJaSipQmwVhb5cKTPbucKvRgjRS7KJ4MK8FE/i
LY7oVd1OR8a1ZT337C7z0c5E0Mqmb+uoe2v17Uvubv/QlhtjaZ2rWZjd16Fl7W5i
r+ovNrc/dzAAUrRiShrU+dxB5pvNUMk8hRWQ3WRvk157w17kPGGAUQdGzHYgW39N
MQj7r1t7qmFenmlpPaS4c2iSrVSr+2LYuwJU/jLJp+4OGUE3jipYYTqhiv5HC1RI
BvoYcAkozsOicJONvM7hr/t8Tt1oq7irwgfBmnFtFCWB0o5zZ62q9Xe8Xi9TcHS2
hnZO49SDiAF11y4K4BONF4WBtxobKTaiMvONKitk2p1bkgR/kI6DBRipANmdOclt
eKjYYDsfFheDa/s/LIPUiDXRMCQ21E9SZyH6+YAJRdp191ta9JJd/WYLeh1sU48l
zNjCsnqaygXypRscuOrk1f0RR14IMSEu57fwpMgP4bXOwNPMt4Fw8XlFuD2Svepu
UKh0w/Y3ZqmOxF2zLB0SZ/kDA7a0uQONHXzV4Ob9bo831Ka3unsHwmaQD5Ebz2V0
HJDQJoqcXOCVHfKzM4J1AZhSXkCQ4dPNCAf4KepJyn7RSZGjHyRyai4dxkP9DYQO
zH1sRRHYDTmpGadxG2MoKpdZzo1DUMhZWJCJ6Yav6CBQ5vWGC3qK6c3HA8EDUYeq
BI4MQd6uLcmnBOhwhang5XTrDhH85PnRFTXI7q5YpgfWZAUg4Vv3Dm2aAVnYo8Nf
Fau1CddXtRpwQi7BDgUCKkgs5aJnJt5exRcAfVs9kS/4N+Z+Nw/F5RzKYT+Y1qf7
c1h2hmq1PqCt6D/ePFCRMYlxfE/HED3DAhNQCwU8nX1rSaQXI752wXo1vxy1Pcd9
WpX7CH9mKLcKH90OpZl+1ryh+W0tIPX0kTaI8CQidK5Zj6MAdmhr+0PFxcvDl32F
/16gXOoy1ZingSFO6GeA4Q4QXejsq0sbq9arrVAz8RwXo7CcMQC8e1D3aL6UrwkD
agwNy9zRRi16H4/gAhSwFyEmMQ8xZRKUFgnve1Mxiwvdko1bEYDL5QzDXvNl6Ao4
wCrRuyyee+fqQRNBca1EhL1JNGMWvMHgspTmdJ12zDbbAiFCRQO5pLJejKlfdpQF
i54++BdVg9VWBJ1FONWCoQCRkhIV27lbbZHFLNEnOfd0e16fq/gSdyiRafCd/WZ2
FgVHPNQ18nnLoK8JeZdGuqE1vsOHMpPiRVLyEskfhjboTGVm1LPOHqsevprbFXWr
dk2pgS8cCpPSRxUvg4KmxNk61qZ5YPn0i7FdOy5P3Vi58hWPdcYMb2Geps2/ReiO
LZ9AKZE/VC23v+KhYFh/EI9t+zgMm9Dfp9wF+OuX11otOknvas9zI8sBm4eaJHjW
oP33lQ5QcCAb1b7/vzzuSmtAsovEHet8y64BDt9SGlTgKB6yzFzgOMOrVtLTgMM8
9gQ+8x54kaxaEn0VBPNBYZHNNavv6xQb2l2H0yEHUnYfnuCq9a12Dnn0tLyFq3wh
56nLFQN5OBJNjee4UQdmBrg+G5Uf6A+v957mZfYeea5x2i8FrryU0QZ2TnNpn9rd
t68VT9vLPXfvDF0NJZUl09dYKi2Vu9LtlEfYvX57WP0R12Wq5dsrkDAtHEVI9bUS
JvCyzbBVg3D0yi0Y0ILX8LhdFzLq6NCn5rtYzLHl9cqFQQHFg9Cj/ohvxrBl0cTT
ZW46GqD0ZJVkAufDRQ0x5p65dcyhoW7uhgRWNQSH3pSY/8s3t28xZMl9AO6EJ7ca
Scw/14gk6J1Soexr6N+St2yxWZaJiK5XN4q0aktS6HGVdayhOGfeshI7xuP0Cd7r
Bcrjx7SJWDG6EZqyu4p+IrLbvnhBpRJrbuJ7jbcoemnnk79l8id2uxvGu56ofs7O
Dg35k27TyC9WF5H0iiU58I6I+e2rKPzpvf1V6axmPYnYi6ODz9e3AaGorOLkxKa4
ADDed1n8ODxY5XThHLJHPTjCa8ae5Ytvf4kgp5zERdumkYEBeuWuj46TyphcQToT
xWqhs4zUIeIk5aTtNOm3Pk8ZfEUqanvGbh4KjZ7JkixAatMTU37c0yT8sm4esVGW
5ekRQBzJp97EMXoD2U79r4uN6AyxBlBl3j5O8EIJ1Yah1iVNmPQmGcHVVQM59NQv
lRoyDeMi6a76dbve05vtM1EfPo9kXWvzW7u2QV2+p501/JIrjRFAaI9/QGKZO6mA
YwYvWiyuTQ6OCE3D+VvBOGvPKjQMGfIoA/OiuddVQ9yRfxCy4HzfsnOX9EvAiz/k
M5tJBcJanaQlSKZprGq8YnLr27wTLIQ8s//tv13XGUNnk+/4dFw09wo277EXrLfd
kR5WxcW176pejCoem0JzTxbCJ1+2i5mMYtlf/mq8Tqeuq0An7C0la7EjHmD7JfdQ
pPvmdHxG3oL/4uIbNB05GHEwjWH8L74xd+AV1RriHS7vHh+tgNAa2/Z5qjHEHZdX
eF/l4VaoAVo3X5OE3PKMW6Kl/kMYq1wNJncOuEJRmeaChoWbgXszYPgThOjOnLzP
wO9LZ7bNmP1ivgxkbszcgqKEDp09m7sOR6lTRExtuxvTZRZ2Ivmm1zUcWsHB0/qv
Y50w7VPsutPGBEcYXlkcJgIhgBYldPchovcO60Q6Fb5cdSnx8OvgrDv77F5tUZP4
baWeMV8rBvbt8MYgBNy130Ii37CuErfEgv5NAmWffMe/iI4MhpvxoQQw2bXxILLQ
dmjn97lCtrbbgizglJmr4B6gUIjoQOleUJk0grdof5RTsrbLqUtafvhZ3/GmXH9V
YM9rFyyPYPZ4q69XFrel4AOIKszaP2cyL7T9NdoxOfwicq2DVcqFs7eHyuWmQS90
D9OiM6fvytl5YElbu0EFJhruGe4EQ1w1nCP+bowKJQ7659SA3zZmKxUAA0rLWitO
J7ahBW34XmjK7VPW5KCg133jYFmN5j/wEDcoUMeh/rJ7Ex14WgZtgyweQcOpwv9p
oBCw8OCUt5GF9ivXxbGqPtc7I8+w+m3BtuBpoRJGylG9Bgtx6J+TcjqNqkCr8mV+
Wd8ZwHGIaG6CigvBrMxyl+jt649JFxjNc4+HvUD7/vnC6mzVOb1/2AGYuvTC0I5p
anxPfDRMvPKX+JhWNi2mdplLbgYIZFOHh5wArQ+aXS/AME17vJEXTR5Kea4EGwoN
XxY1VSUKl3OBXFCId6IMPv3/HOy5SAfxykhtTxi66GXNTn8Y+pw7ayEf3b7Va4+J
UZLkMmQDzcMt+nHKs5rKVVX4fo2wL9PXkOekI0ROUpJJi5x028WoZgRUPXtaUK/1
SIea6bFowwXSR1tngNy6hU9afxCTQSVpLF3O0+gNpAqkfevwcYZmBZF27uLKz4zO
ySZ+Z2RVViKbUuUaA/zUiiOnRHuvRGvwgZ1kCHsmFpc=
`pragma protect end_protected
