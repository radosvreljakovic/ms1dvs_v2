// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
pUlR7x6MnF9Q1Adr+hU6EPK8Zgi8gud7QYg5HWu3bJ3RVv2okm8yvWHBeNB6GE4SU+n/QrNBSv78
1PBU00qk+rQw+7JiljCqQZW15ZTSx9W+c7L9txtx9JJqVkLjCpkNRaWtIAGU+r139mgatKqx3RRo
k/2mlSv0kSaYhZTsMpYdSLdn98p+FLYz07GreY20HuZ2/3TR8fwgORPyDpDRf99/es1PP7WRmhTr
tosMMecxxKHJT1IRoheQT3jBMGes2V4qdt/0o6iHKhKP52c2MewxvFdEpJtFOdjvPruBEHeO2o+f
6zfhOx70p3DWWa3zhnl97zN1Pq/jMyVJSCbk4Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
fq+/0cZ+2g00vIcyv8kSglMLUURIGN2cE6xTfVUnazeY5VSIu4F0508gEEDadWg1uIsyfS5jK/iK
ZSstOiRH98QfICEIwhmnkhMdFGnqruVWn+hR/TR/BDX01GbPo1gCFb9RIdlvdbjjkVoT3gg+uKRU
w+rQ3dkSch1ErsUQ7imGAbwbfQ9cH/JS0vj5z9QDh2HDKwKjdNd28bzclr0rEGcUSYQ+cQiqoP7D
+kxOZqzyYQlLGme34qxxgrDqXAIfqHZ7MtleasL2w5FlSHHGwlc9f+eAyI1dDzpYd1PPKpyLW2C9
5VVVZugKOj5MAvF97koAlNUqlJ7SHYIEXppn0hz38M1tNOGVGPN20O/YMBIrY5abYDJoaoGjAAey
JVxeT+caURjoKlpGTK0nQTrg5Vm1D89RNKqRl/fLX/703sGLDY7OjPRU6r5PBk1hhauC/xtt/CcL
dBcSCMCv728LnF6dZS1v1hHBXoLtRY/IGPZwTMA0seyqScKWDYsryx87uIQfAltr8NowEHEQYnoI
i0v3DuFx8t5QYiSW17kAQvebiBjr8fivAEfEzcajarRH1o9Sv8lZjDEfqcKPjW+97cOv08en8Ro/
EeSPOn2sAF7M9HjwMF0K3LHJ8YVJ7oggxYGRwjrbwpzypnDAtw9G5GmX7SU8/kG1SPlc8PmAUhKa
gFy/RV5n+5a7HvML360qn/FhJVWBKaG9jNDmdIo1F8KRgiMhe6eIROyuy55KB69s48W1oNUIQZa0
oqyqV0klaZwhHmzGFpnSMYch64a5XzAr1oAh4r0OV7Tlvh5mnQgii1JobdJmuEblg8MljETvYCpk
8cHLKaiHL8+LqauIHDRgmwKoixwIa7hWKioT3DfPRdXL5hWvv4f1KZrDaJXhshFbJW+H4l/aGIUl
RKChtcf7IZovdrkzO80hH9m0nx1U6BqTmFgJsr0yOmLUaTiW7yTr8/eAOWDyqN39lbX31h6110nO
LcLG6IbBlbuzVlsUb9AI9TU1PNRocNK2pSBbh30gdDXjYfpBPMKSkNSP4/4auGZTvzvuFizzJq7Q
o6UMvMr0BueCstJihAvnQmn3UKYoGxlAKkIDm3c0mZsfv/JyS3SWwytdNQ4RJPo/u3AONrZWPOCo
J0lvPilEic4Ayjk2YxAculMrYbyIRnP1GD9anz0e0/dj31PP/wTYUtY1ctAhKUXMEhPMjblku4wH
xdetExjsE3/Z4GCtA8skByK2qrst4wwpGR2xsIRjWitPYnutdgyOP9pAS89jaK1yQBkm4mQWYHwQ
gBJuyyDmYBInk7vBnxbvHOElxVPa//QeG8hwMddG6J0qcAwLcqrH3ser8PpTziw7aYAdvGMyDQB6
5bfYizmHchtFK2ZaXjtIrfs3oUeahNkuJKEZQuGv7nodqYu3ppHObT423gW8yMt+RSxhTA4hBZaO
z0WH6vLz+dJjmF4m+R7WJvnQpS3x0rRfx90Pj2e+Fjtvdl/+3VM2zwLmAofhDKcmbaDg0lIvIGww
clPJzkdnPF0/13Y5vJzB14UJ8qxhhgv9mlSam1jVz+1g39z63sCucymzgJudtAmg3WCILwtnERpB
EtNsKeF6gbXdnAIUQwZbJKVIqgR/KcJ11anOrfbjXWCvnL2r4mlB/rFWSGwzuO6kXGBBg0s7ShFX
l84EnuoRyI264g0la7zvt3aZrmaRh9QpdBgXhSI8Sg0xHwaaI7po1UskKFwnm1szhXUNsbExpOf1
Bqvl1JJL9QCxD7rPCTjLD0+fOjCCNyRR49NdB2J/gay2mRSLlto/0sH1NkoL2oePByFMQZcEnVSq
NZ01MS6MfwpkPNCcZmnutsnraL1aVmb204yRRoxWhr2gdjo0GcOVqs3xtpHRhC6uCR38PSoUsvQO
9qs7rY8NlZBU6UR/O+S0g2nL6YkO8KUZtBDDtBnqXVcy+52QOBBjRX3EJoMFljpyDPXU6XHqnUu0
01cy1gbdTwVEufePwqtXZvGanCRVIeiO835dmbgWPhschM0yWQ4xTgwwiQTMwAXcEc0TsooW1zMe
2D2nVzvK/vuOGOGszvKaDsch9Bx1/xCgX0IY61HKW20UTe6JReTMC3/Z3etHCYmS/MkmTnFZwNoK
APBY9opjCIVULE6ee4bJ+xfbaYUNFRGvzZ80JZI71eHeSD7SeJ8wE/xLvbEcNn+o3QGwKX2YTm8H
DKTzIiqIGnhfoIy8+RMvEXT+yyUvQ6N0B4WcpXN2JXnK4+LFOeB6peoIF7Ny4bKMVZ8czVTAeCFr
+qSoITsA+99xqqoqydyypyl7aaM1Uf4eSXKeMa7r/NMaxixu/MGDK7OtzcYmteBgDQ3d9IWNzKGf
ex2B2Sw30G/XJ91fTM+la/gmsgyYLcGP/8KbjfLTFUZS2CDSah7+0xn/qEL108Z/CE+J4R1oFXuf
4h3QA72lz41MDE0X5Dp5f/878KajvMZxCDFtQBedr6Y4+aHmsEVnb6C1KAEQF++bYd/2XkRj4KG7
9osgyp43n1xfk53xLoUMewJVe2IoZ68kKIczbk+m5uQA3KKHtVT/BSiYw817t8HxXJ1QLXCVTuCa
v2d1o30hdr8mEFk3z6VokwCO9rZoAEgSkAMZfewfhhQMvXDjhM8oZVf/QaOlLR4wWptmyNvf2Heb
A/0ClI8CO4wEzDUNXsMY99Xy4BJG5IRBcTTQ/bnyQZp2+7xt8yEEnTeY8gZzFas/+t+Xe0jA8NdY
ZGJN9hz42fBE1DiSVdRzA0/HjCc2F2HGN/nNkASXTjRMTh/N3RdBsiV5di+QfCypYuR4ad3s+9dS
D8XuMcGAIfe3ykyeJKaYP9HmNiPi/YATlh/u0OyD7V9X+omZEL9Bwf6XTIidtk76MYgzjHJHFvNE
CTmKqR2MIY7CngKoiN9m5A4Y+/Lyx/CkcJ78Yuj7gYj5NOcE2HRHj3tZzvBWpK1/CNt7SwZ0fCSp
YW26VShBYOWslVc5tyUnyWAMq4F+hrBuyjnPqErSbOuauTYuoWaK024cQoIVjf+FtCnzSMQL7HQm
tTHjVRGVCeRhCdGPmvkFnetu2fgqdB+keHgffCq2/nYXqyi4t1IS4VtdBJ00na7bdL2SLcTFQUlJ
p6P3N74sTnf2YTAouFmovqTeiqW9hvG+qoEK8Nc6kycjogowxiJ8wFHLNRA0ZpNLdz81WjyRv28V
3kxHhg0AJW0wHCuksKFtgqOvQvOz5N1t9uxlSQo3gu66dHpUh+yOQ2nR4x1LbFFOUolFwoXu58+e
+xK20aDPezp6QdbkLw+Ib3Bu2AAog3cK8r5fo/4vPWmeWRvoi9AlDqzuZ5ifyp5U7Mh6u3pbdCdp
EHFn7x6aYwxIF2PNhO9MjGpyxRum3S8AgzRQuHT8ufA5+QaElBd4k+qGwxo1r/Gt7UkyK63FgXim
FqV7Pwsc/a20hp59EqwTH3dArqxcCn3aJ7sn6UAqBj6uyqaIdexaq6smAFmJmEmHm+aO9qsU3ip5
PYBHJ3LJCyps5qphlJigsTjqBUe3AD1UaG6+Xsvcpmt9EDFRmZGLqxr9aVRa+gWuh66peSIypRnF
ipKjVH5E3IUl2Ddp2L7rYaNSfZdJt3FzK1DUQwW7XQ96USh8i4aPFSrkkr+454SZk2a4YEC6yS7N
craSZatXpQ0m8nC1Tcurj7+0wNi+aGKzMQhf4/HXcf7/1N65FUknndnUpFmhQqzxY5eThehvSsq3
7Lfb4CglpzFLneBDeiClCbLq1/KErmNajZTjuPfwl364D4Zaa36zLc7xz0ZsbIF1gE7eJZ+LWb4v
9iM1Xg9AsIGnalTvsT1+irtyk82T1ATwqct7yP4apIVT+dDa9/uzf+PTXVTDCDc3t9p/HqY4LUkz
iaW+3aV2eujvOoNodwpIU4GeVNDFUf84OFoJwDVfG3mEbV3sg8y8bfH92j1aIeFR7werCI8ClwMZ
B/s55WH6sgbnMfXYFj+1kvGuR75V15VBMYubwhtLWh3NGp9v4tDMePvfijcWUrDf5fsaaFcAXBTe
nnB7gDA0RXalEvy64VQe2Dp0KKZTz45MJW0cQ6mpb9WPKZVm8D0qeaVokr3xcjIqicVjZ1w/vxQ6
dLcP80bErEjeAESA73XtAEia5rGjd4xZUAR1FUJPQ6uy77ogOThTf3sTnhwtRmwTuDWczCrlV+IZ
JhxBOVElSbiB/bhHEfk/WMmfKD0DTNTXGQeqmRZYPVGCNMvem6vO6o2gP0pktKn7R+iYXTX8Drq2
bNnIfvXrILm8wNgvtdC23ykYAGvdZGBewogYakLJgvcX6FQAWByyEOB4wVtG/zTxLhGXd6LHRhnH
yU1WupM7/s+6d2qJe99uB/Ny3g5lNV2XV6zk0aAbBgldXLLRWp8DCVaRhPQXU3aqfYPM1DOE1pyn
1UKgEmXHLVB/i1aGkEBGEt9g1wMQY5QKcWSCLKi28vJ3zsMIsnQn5pKctAHe4Qs2tVi8o+Qc3Erl
hcI8sdePMLxjopT5BuqL065TlUICf6CC6rUAhXBWcFpfn4IZRXk0DVL+inMMO7W234JMFnECtojX
sRPDlLvtjbt8110EKFKGdgqelE2/8/cE8I+ud0ZYi0hb8ZNlIYPUCNjcGNoL/GPa4+JDTxv5JPi0
w0zrMUJPI3MbfYrkWxa2pmMxdU07J+D9XZK34T4oi39r92kAhJlduGNavFaDZYOo8y1EYuSTAQOM
JDhAe6uxGlGr75Fjjgr5wEZCcvDQy7x+pDNy2/FIrv3950Cfhne0dU1c9/szIzVfISnEJeqa44Uq
uwd/webvnl5mJa0gSV9JiSkl9TRf+uw4mKHxaU/DH+5GFY/ZTUUWyuWl/kmDtFh+DnMvcTWzODXX
ssMxJj/Qrx/XkbWocD1yVLqY6vBw/GFehAkW7IEm/Nc9bqzH5algB680V1qXYxenkKl/6j4dEgC6
Tkj4WXt0M+wxyFcBFjUF6Y92xk5OtApH40nxP3QiatjdOafqVD9QwJI3kga6KGe41C+Tid2Cc2e3
/i0Cam2TdTI0gTZ30jQYOL/dFLFTGiWvaGIMlmfr7TvWwXtx4EVFN7uuZnTpF9COTyO8UN/IcBms
SqJK1AtfmOmeksSGfErknBL/bazgrIV68ymp80uifiz+KIgxBMIyw/OdeVcg2aUAZ3ORp6lnRCEl
IzH5Q8u1m0HRheVFNqMv/b0FZhqwYE3fllmasMeQO6YaOlXzyxuEZb8h7RJvCSteyBgdAElSnEHo
Th5xMtAailAnRq6YAVy2cMc//siugr7UtXrhgITSqX4eKMbQ7yCf62MVcr9dfhe81+Y89XaFSAxK
NcMnzcBrWMvC6W2l229BmVK8NYOSH8AlxVpxthc/ECyci+bu5ga4ev0/QiIX+5tN+qkLaKQMEPSB
MCGjl3dc3oBSoG2msze32Pbmlvu4VIgXn5iuVq/2ThvpK/nxCOR1CknLRvEozsIlMddKN53KzbLp
X3noJC7eWmqCV2Bv534v8E+0djMS70jme0onpbZC/Ux11vBsAbvFXttAXh7/vzqmjyXUnpm7serr
29wfX4GNEsw09d6BwcrNNStKN6F2qBS42JYIIz7neTaPMfl4sP1xFGmzlkOcmc3iUEW7Bm+LVIZa
9v8a/xe/Ih3uLjC68ufYJafXxX/SGiEmn4FyarLg/TCN5bavKGzZLVFBQdH1YAIzLWY6BFoyno7Q
sNLXW31aIBMeF0hiqCS+1xq8vZMcD8LtdWRWWuCmXjpdan9sZsB1OH5f4oMhME+jTiMzIzAdro3G
oQlQcmraufC6pAAR5jlOvhu3X7ka4xNAQGxC5vlcqd0ZGINu23NEEERjdSLX1qfpEZAX1argUstM
EvVC4UPSE8xms8BY0P9evSaeowlPrJtQJgUzbRPga4UaxhPUJc+6JL+mVcocs3qsQgRrqctVPDnl
aHn3y8R2OerBRbUHbXGT4X5NFQdFx7jQ56nwJJXpyIV89i6ycJ0zKCU2aE1IPJlgj0qm/xdI3cxh
BYxH3MSs1AnpyGpUUNEV9XkdH5tTzsEpryHqJ7YlQgYVa3Yc5KygjeUrULgZtEAXE5r4d43RzFQV
WTRlyJpAluXIpi4ijzgx+nx4hcngoKv5O7TBq4e7Vbm22tY8vhd8iJpnWahVaXv3YTRqXzZ75Pxz
WfeulQu0/W3xhmplPRrgtBA6w5kKjiuROmo34H23c128alrs2gMYcZOMe1lyq3pndzOFQH9Opf3r
ryml12mldvWx5hdPhSvzZ+NJkvQ/VxaOcxH4XJp+BjJ1woi5nVUH2n6Cv7MDdPVU5lW3CM9NTvpz
v66cXMGCN5LFn13sB7R2kL9kV5rwJxiune/y/2MfcoozupBFzb+PJ1LTq13W48PHVZv7/Jk8IihL
MWsYMo+y11aWsc5yvCM7t6k+TgUXwqeUnODTQwSHWSyt/mlTmEcwk9+Ql/0j8ovA0kLkJdyKf27L
5AburMYDC93fdZusL/Vxt3TL/Qscw1jHSiFVVolX2LfLBKZg2Euo96KGZUl2q0IaI0vA6D8k+XWU
P0gViJPp5c/h8xuwxMnnfxcQYy22LhoIPdTObIqagIQzmNel7L1hzTUDGHQlnWx+jdPFk6/zSInG
j8WhH1jv7AduU8aXp3T4ovM2k+qVGVMY3zuIayNcfyoKVzRTs2DvWgGOQc8vCtgN2HEhO1RIBtDj
TDmof/vAlBCPjemptzBPY6tNXi2Aiq1oQioJhNXe5+vf9Jvsal925SSdyWt3xkzTl02My4+kC4pg
NlE5zAUIcO5JjfwRyZNx1snsylbd/gNwgR+QS/Vu5EnIv+5YYesmNuPOQ5upMSD4ckB5KqADRkJJ
SUh8se+WPEalJoNiuJwo1fvT6WPxeWMzrqH51ZbdGG5mWlCUYmRnBY7zypLNolYCxjn68dcaf+qp
ykDmoxE1cxe/sAgQo3xkwGrZ7TjtI9VPHZM4YY0oSmMUGdNEtuyoqF1P7gfFSc0gzwB7GuvmJ3UT
WWD1RH7yWBntzJmrkF4aaY1nb2yZDiiEFDRgHRwP65nWFdsWSg4ketUF/y2ALPifauxGscDiez0K
6GkpnvdVZHLgMbn4/EavXvpkZM1fA2wx26dl7zNIVaCgmyNfAY59hcwh1TmT6fJ3BgTNE35B+RHE
sNKYGhuCQVnulNW8sh/s+iQEbuFKlEPmODX6G9MFxwVR4nJ7sw5P3n+qzgB4s4tKsQBIFbfwyQhC
mQR4mgQqV1bf/3mlPICl92znRfqxUz9ZCTaeJqjcW8838VkQ4j5JAr8Zde6BU7xR6lMdJKDnwwn7
VeY/0wd9DVRhk0wUyiS+i5v/0mTbUNb9eZ/960bbWcdYRVamqgCRBZFIdP178Kgt6rXn+lH4K3NJ
RhEAEdhCozghMkFGYecPMX4SopOLNFkQ+d7x59Gy6TJSAikb2v3knK7z9EthAxr8DLAFwZ9MuHnp
SCA5c42+JlaQKkHeTWN/LT1qDOXwAF04W4L1Y6KMLCIlWcJswMpp7yKdO3w0cMyUMLKajhcwBqLJ
YpTP3awsWEvFH7KMgBWhRDmA6RE5lIn99vhqmwTiK2HGl1VpfNMsw/8uQD8AG3+H1BVGboKL65fW
2MKSAeff3E50CiHjOr8FDE/TMtWQOjWKrbOGG3MDLZnoBzX78+nY2uXIuoI/aQTX1UFl0XCc0u4r
Ko6CexTkUxHyS/XzepnJ72rHcvb8fuE2PYnEQSepGLQSNkreBiG8oU50aKV1AtbH5MwDfGiT6gVY
oARpOhLrKeaH7bilIltRA5AbRohPOfMMCul3cCJxefAg+TC3Nu+P3tzviDURL6T97z5fglZ9yr0u
0MZ0g+n8pcAKYWvCQK/iHZ7mKU8Zud4VGnIJVfVXmNI8r45PwvQ+BIqo1R+XC2DbiVSZgTykd6Ee
jVoy5Qa1Ab09hOYjVcv2Xkqr0jfU4pswZN0fqjs6YBrrrQtxJhyn2LJctlt3ym3rM67mANU+bSoH
pNEn7CWDVkc4TDknpTRL40kf8UKD+sgaocBH432yZwRVUGCvXGx1Rn/f9HjHN9XHjEgupMKU/awo
kZ8GxzeXgxOxaDoZUYmpABOiCFyOkXwUf3jbJuoEAr8C+T0EyXOGx6bDLdesqSp3BIV0fL4WkPIZ
fxeNhXFNj2WQJp36pnhY9ZYg4GsqIXomxxUz72oMtwCZD+sHzqXFp3dpSD8caGbsaNyAk7o78AgE
30X3V2jIq2/Xsh38i5pLDivBRrDvdZhhpe9OqY1lhSei+CZ0nmTmeuFhsucN7fgVW/5wE3kKaV7t
WOmkVqcSApAbsuJ8HTyCvsSqYwIDLLN6KMWcWCLxR4G/fP68EYV51ZVt8+IUc1Byw+PdFTabcsGS
+O5PX4Z70hMNyHRN0dmtokoaVMkgj9ku0pzib8AL/e7btoE9gozSejV9NQEeiS50jLLGoPzKLbbE
CqPzz6O/JJ6XED+xoPBsbwLiAtKIkX/DKxZNOevAPllUolR/PwT6adNRL8LzgOEi0BnfuOuBUjkd
SoCLOZq/Z7ez84Q9B+dg4RU4BWBfubg9AFEpALNBJFk/r8RTpu4rFoaNGsFaS0+4JJhebfNgjsrB
tnOuuuYp00WjFgbk5q9c2jPxZZaGQVS9kvrCUOY9iO/KiUu/BZQXD0eCCTtoN9EYsLtFViO8g33o
Uw3mSdfnFrzGP9X8Mvb6+Y8kyK7lHQ740GhTvl8UMu3Ld0I3P3A4YCBwHUtNqhjKkV+obh9HLXbQ
W3F1s5zLP/ltUZoGjVBFC2tPCUWqvTGp/e07sXef4uW6XhHKm3kOw599Rtd0LSm8Sj/RmjgOrQhj
ogeCZVY/U9lzeQdJFp9q22vC8bml1juuTLBLTzPIHSONeNR4ZdAOmn6D/V9uJUrvdnqbE1AMeERu
vbkE8aaeeV7jlpojA0mPQnnrpGEwFzAQPqa3/8PcBu0khqvchAnwEbvolknAu1QHyDLjRBM8A+Rc
CJSw6u2mgHuZL7dCOHvYA8Ao5T3XErsILOuuGQ0yjWK4WXH8JF8hViAAOu1wZOPcGsP+M7mQtYwV
liI9pTYpT3typsB4hQ5zdxpv+PLKgo/zaRxWWNCbykYJepLqWRaHk1Rs2yDqcO0LFGbxTc5we8G+
DADlppo4NMjLZnCkrX3HPhnJ/LmoZxyhxjlWyJ5OOgoJhNsgulQZNwxwEPbMJhPOUCI24s9NpEdC
LRN/ZV/pmZB0bqe5CWVr559IKW+Og97ajSGKqay+LNlY1XUtUyFtSwAZ5jG1biK5W8imM6CJtylu
JIWnFyTUwlhG5FNhDzv4l+7s9WXOYRFhI1fepNe4kKFTimb+pWGT6+etXF4JA6gWfkRI/Zfa8qW5
13xi/KJavSkVfdIHmIlH8/8QzP4HUf9BtbmFXXxdy01B+yu4tA84yT5UJg0z4t0Pf1r9KgLiZ5/0
5e6uspYsonxIRUGEwK0YCzdsD+qdnlPS4MPqggXZY7USof4hx4+MpNLWoK+sOe93csaGewD5BNVF
MQHdFGG/y/8b+AKJCu8kDpeHeiFcjxaz7ZLWxYq0sSFXizXtn43ugapOVXt5Duv6LchNmWbO2Vl7
n+BOTYZlXo5StvpuyQFDBV29tB1RdQ/XWQbAKNVsXXjI4RDCxpVyH/bJtV9rW6t2wbRt/qsg3fqf
xglaOaS5gBAHVw3AF9EVrzyh1HzXPUHhD+i4C1bzcjPVOt2FB9lmD79RxG1BAQOcu2WjqxfY3fKE
ZyNgJR0Efftcbp/Zpf7bYmSlW4kL7z6hsGV8w1HF2joQRjGOe8yUITylMBwNm1FP1bs56ehuOk6r
IznUyE5Lcv6INu9/tVDtsrMvOnAltBqBqkHf6ueq9zHc96bjHLvmSVT6lki2wDI6PKeS0AFjbBdy
I+6nBoiRg+Ax+xi2+orV19kevkj6pjcgD641PCtdKordTSAOG8/rPBIA5hXlEQHP6IMbbt21TmxL
y4aGzskduz/MKiEn+aToQ+fGhwtEKUZd5ZnW/hqdtRpdi6CfiG0EuXHX1K4MYR3HTwtXOjuMGQgC
5UhPCUpqwUIFR3bYCxlyZVlmPMvu62M5ydDJZjD23vlUIyjWlTPgbp430KoJn+qzktfUsJZOMyMt
yLowotU01LC4a2pM25XSi0OLXJpXczjqOHNW8xJbIF0HJ0yHlsD2ndSqgusS2F+0DYtK0EKcitbg
aYpyXCbj6nHeARnUkdF1c4WcSEp874DoYa+rZqkakIgg6ZGhSB+sVb/w7gjbwxnrQm7Vf7opFxbi
vQRG6b1/CXgHznUipCu5A9lwCg2pW4Da2yrP1fP0/J6qtlCw+3BF7gEtLjC8Q/bwlfdpTcbl6rjy
PXf6XuufnChLIjIxroqFQy1N+q+kS2hZyTiEYJNX4tD0BDYvz8TWMTg7Tj1JRw1yQ3vpF6H9J/t4
J7dLkpnEibdyUhG651uMmTxvPHiuUQqYL48qqJlgsiOXr7bCF7doE4I7NwDcKB6dBKG9fI9lJaRU
2C5W5etwtucIkJpGlz1H7qai36IVcZgA+0V3PYb5ylaNXVM5KJrCe4JLD4yzBoezdQFsBZyz/VVS
lRVwxMFP93DnkCVoWVpjBrstijU0lxGymFcM7YEukvcFfSB5sHPmbr07IfP1JPGFxd7vIs7fOw2U
x4e5Rg5zOCWQnMAkw2qvbG1jBGVRCF8RJoodKXjHq08CmF/FHFYvMLgXKgsu7uZlJpDdlCMGUAmg
A8tsRwXdZ4oMzOVCzd5Kl6M/a8Vin902uXUeiPQS93IpkFPBuVdRNk0SeyP3uTqeIHsX2gNcgs6j
XhGnNE4plghs/2IAg6xqqrcUrUuJuoXw0OwnYLevQv/xmxkc2con4s5tqhZBJtgRFYoY4rTQUO+q
yRh54Zk6ukfDd7w4ilXvYCZ+IoJJqJXeSEyC02jDbogtPcZo6udadm2cmtILwtImJIPOcDFCzp9d
j/iDs8OkTG1iLLDVVlLR92bAxNqYv4pZFek6KTViU68OYTWszVpXvaaHYIJKoMuFYkXDsiLeIVJE
y2t8LrsqrnQY3oce/pmolHL7iMj8A/Z4LdCQ2az1+OsTZxcwLtN2PS97ni1W9wVqr44iR3I8BBy8
K56DCuRdN36PO0as1EcuGb/R6McififoWfSVX3eR4NesT0XKJiSEtrjoF03aGQy3S/sx8iFaAI+M
KsuxwHuhDDvJSTwuNmXbLexOuP6MMVwVJdjTFDhZz9AlEEWfU48KXVg6nUwOLyUaSZtHpqYYOUsu
yGrSxU3tTTH9/Gh2NxSUeUn9ZRhYby0RXCZx25SryRqWairQrBZ3AIzS2Ycet3/BqgV4/9sXDsE+
CHS8K3TDaMZOIIDyF6+5UZK7RLd7qFPc52mMoGJEZ0HmhrglEemPl41GgpBlX2fPAgvUAZjo+Eis
kDsY9warQK4COGzc2SykF7INiXD6nfz6h66BUvuVFMh1UHh5goadUbn8OJo1CWVNHwOVQLHyAXSg
HVIXdEDsS9MRqAsffHezbG9mSy5EadXL2Yjb3lLly+07YNONzWnZbToycaVxcM7z5RganKS7qZB5
mnirm9f7l3oxywce78irz9CdOsfX7vXVidjoAZ+D5pEYq4MmFf2K+om+hcBUNpXUFz5y2FUP3hl8
lA1p+xRlHebF1AXIVLztISBorb4W2XuBvluVJ4y6V06JNXtd+LqQrlSSTA6zT+LnGRlHEi9D4f+J
rmFvhVQaMpSnHHBZuOVeQwUJUt2bc1b7rPj5UKLFZu6V19PZQfElx24XFtDM4EN9gVHcGV5/Y4A8
wFCmA4oH5vl2ZErkxzgHDfH4GQXsQNG4bVPYiNFPwiGDwCL0L6BCtEHiD5Is4I36BnzAH2otpqK8
dRMbq/SAD1WlYGsELaNHxuMPBPf61j0NJ/XKvhD0gWpvj5FcxAd8Q60ahCFKCPf233wMykMKHJ2i
6MIF3CtSDzYOsmkQDkvmbCkM+6pu93cFfKmuf1PKgQfVxxXW3cTdDxObn/N5NuhrKgLEjvOXBU2n
boZGpE3xha4lnl4Tbh4v7z7vgDfA7fY4Jia1ZFoaUYlDmTYs+yo3QskGb2c2Vs5LnDK9ctFRHRaA
UqPSbrB8IM1DgFcsYMz0RciDlTMdKVgM+lemMZhgrSiYfVOn77SkBnLU5jltIwjo6Ur10Ww3i6Zw
e5wHlqc55WX+kJ40gzNAA74LlXGvl04Dpe2DHXGcd/JisOZYko72eE2q+ME5mYPHGNVl7/C7d+4R
BfcnTc44VBpx+mcQS9eF89PTDHYDC5McghOWXQsD9qW86dVMXJgIfjDrNuvbwm3izD9cl6IFLcqr
D2DYVv6rlU+ClIi7cwKp/2iqv4VqWLgac/Y8b+/BBZaCUJVLfeV0DZE2XytlHBJMLNk2+Zc2nNFH
gLLvHzCdhKXq3SZW4xxZNjbLYHE0YUK20b1OoXGfT4EJK7xUk9hmMLo4/2pX/An+sGUltJ+Fbt/E
kpAWD3CCyVZGQ7VIe4pJxKSiYkwV100ZT6WKFCR7LnmZPK9B4VhB9rSmrXcVauVz1DTRLaM+vPlE
OpCwW4ko2hs6SpMLhH0zzUCoSFo8O5Uahdhrz2He5SMTDq/df3NbtgTXVtvoLwwXMKfzCmaOMCRJ
8OYVw1iVAaLurglZGPYq6bNymjTO7Thpr8hLtTmk6ZBSwCDKKQvQxgcwmdejr0y7z8tF1aaj99KH
amJKtB33jcjfxTV0+XQpMOX2cYO66l03lZxbZv/phNgXOuWxIVNkcsjMFuF7FdZVb4J7r51OhmxI
hzvM/tGe9DvXlmBFLaUkE2/1+PRHZEIfzSiCZbWlUfAkSUbgVOA+pDvPc5zCM32KlAfoB+ylCB69
y1hcMFFDiwRNtAppSKVWvmCRhgSBchb+KjQLYHvWkGi51jncnxhOlZolhqMEY5yw6bq7Ka2uVqnV
aSnjsA3eIoliHFrhHKioQ+E3cypA5ym6u3C3QCisj9Nic2BdxAUlbj1YJV971tSku6B7U/wOIufA
m/+uahfpzNJY5I4Wm+hOFjkaLPLcgvTNIsbcdYcWiXfZoVGPjbM/X87awuKmSDOZu1+CPoS9vnS3
JZ09Ca6XbyLyANAZaQsoe75Z7CMOIkM4wDOBe/GYmPWpjzU6wrkfXoB+m494X2eGVyvW0bgICuks
3F/y+Ns591WBmszISEkpyjEz462JZAUQSGqvwuhL2p/Q3bgFQGfGVRnC1MkjinbBtljR39fqEiMZ
/eWoNViVm2+OCRv68tcKaAq/2M/FijjJe1ZCIxBgbGl+C0uvxEmNM/fkvSkCtwS5NeKfByoTU8Q5
SYc98MkhVpE6KuLcvd+4STjTKouaqdfmDNlxXQxc4sC7AD1+GTqHWgP0B9+VHR75ZAynsvxOSSac
XrFcxrDl03JzBwlhvFGEwKh57dBj0OivKgePmv9FwyyH/Zpr3iQcwHI96emusEkrPfcdcNoeAH/y
gdGLkcp4pPMo7geEvV7sEubgr0G/PovydxNr1Tdy31y9MbSmeFUOQXqB93HI3B4UPDUiIiWP4UFS
4/KNp3DtOk8bMTQN2i5upLziJ/2qfdw+tgnYMFLGo7BilwLv/C0W5jrn3Y58FwEgm/Mdi3uDJu2l
DGSKxCSUcrW2Cx1H3Ey2GrPY4yrKrhj46TBVSnJKEE7DoMJSHhdgbMwBvN4/PyPCLW3X8KHefihR
ox8y9+gc+WvkUyF+z3GI+iQUIZFjvLMr57xCjry9M7oe1YjT6qBZ/AoFA3lnW9Xbehws6eRRPeeo
lYflkntBpSoNsu+nbhf8vW53K0sNTJoqkqAloLQkiAVUM5LcShSDpXJ3D11T3tlt0p+EUdrkY5A2
SjWiXVzczEU8OI83Yg4IWac6qtBc5+/eIAWJ7+grcJwAgeS/O1+onOcGqWWA8h4BN07CdRz/1QyS
U9IfZd/s22hkbb6iPJt+YgDfoVNnRYfLKDyQDFfM4wj/f7Bdaix9lu8aUmZQ4voDNEjdj5l9pCK8
gcMo7ytSW5HJ4MwJsFcjoda0Z65vVrbS8586a7RJ97TiXw5Yor43YiYeUG3mnVIE0Me4bb90poQm
K98SulmFMkiZpfsuzfhXzHS1nRVD5DAyA+kJ28SvstmS6ougYa/LWntHMRxRZ1F9H5mEbn8/yAtv
h4xN0dU8YeIDP8tuGgWGfpNsbGZ2UfyWunB2Hpft7VdITL70eLvqnCYZgWq6Il2g+K2pNHzCGOqd
7IH3cLyBlbIjwfQ1dH8CGGNt8B3mZqRAYumlr1zm/BdQZnPTrdvHwlAsQZwkCjGAHsyCGDkEx/F2
W3KNO/jhur5aJn3bu3ucf2bFc0gAKBOgK0DdnAtIy1hzBc9Zma8TG+IR4HIuF9cbBcnux+0XN96E
J3sV8+12vxzU9CEB3K9e05Gsc8j6Vrj5r/HNkRsWWz5OhB5KBMYc8J+xXE+JC3JrYvPdmwnYIcVi
sT3u7J7fI4eBqwSmrAYPlIbsRlypbPbNjFI9VAHsb0nKJoRztE5JkykfvRLAvonFnRzMX1sr7R84
sUikohdEYM9EdTGXgbrSBweUEr8pjRYx9e/ss9+Y12jDVNyy5auUtjqiX1mQCGx8C+xtYWU5n6CR
EIQexG1vfvEIZSSuRI5V8OfWdnFy+HNCTqZDmv4B8e5rgM3h7fLiNwYEvNRqPJfB+WN9cG4Dg2lV
YOwif1jwngVrXoy1f51S6ZJY0qeoSIQB7MVHz8ZzxhC0j0X9NGlNul94VBmxMJB/kQTVPsonEzod
I9FCAiV5j/iRVauBKZY/kyFeqnCCkTzG/Nh90qTYgC/JYF7BTUDVzVsM8erj/ZKjzxB9IkcVhAHg
sO+zgUnBPN9x0MBHG0F5FU5ENKaUpBpHgn6e46ST4ljCJEUeAleazvMPS6NAxyCn35ubimrN1Z6P
Qn3B2AKGlsBlCz6O63gyGZ5/jvvRrkketFOwPE3un+8u1Rrm5OmzkDWmPUVqprjwBIDC+V/Rgq5j
82MJcqaPSCa4GsUfod2+jKn2sWH0AbU9QUUsIx5mAK0Ojl6WWgLs83nsh4J0VYhU2P7MKQ+apGuK
vDSh7Mx3dj88QkK2mvDZXNIb7yVnEyNLDL1RDFuTaliD20kRd2kliTi09dcbpBkxXk7tfF2kPvmP
7cy70GayYkeBUSaIL9bYlZiElSEj7Y513VpYnRu2k4PcOsSEVA/ZrAyPRhdo0Pp2qaTRBBDIxmni
DAIiLv9p1HyqLbsoeEV+AS+2dBDajyWIPgJ/rZaWTX9qHtTE7NjtnoxNos9mnQUJg7cDYAlqeCp+
MdA4Q/BGQbc9bvjh9lA/3uF5tq/WaJtjwd0AbnOeDXT6ZBdTbe9q+HvLpWyv3Kb2VABQTWmoEtuF
81zd0CFXF8iJJRPwcpOJqi7q0krUhxRIec2atwx9BgR+eoPWY6HM+VymfDdAIVHR37gCq0eXezKP
/fEe3HLoz3UwITxmvTEu99zgos5AN2gAWiee1Gp2t/NpA9N0cnXqlaqKVWd5Ip4dvNOmtFdKdMFd
4Ihi9SOW6C2fSdrQWdLAqHUvFckwjV5IJoEJhfmvLE877WFOThuOEi4PqutntafywY8DqecHwf47
4RkXu8MS16aKa/f6iZ2RP/uLH8/BGCuUQDmLYXXAWmWEKy1xYi6CCgok5nNbRBp0dgIoXSFFJArm
FwuiIroKsxjfB+jdBE1j5h96Sn9tsIXZgDTPene6xcFKRkI0DivOEMekO+cUcDhEvypslDYKy81B
wh3ywVng8QDeGi5P1NKjYsT0kwA3lakIHZKq+6xM1wfoxxZMMtU1Uhf+DWpBD9Cnf4PwbwDqAUkf
HJ+gBVm52QDQe+093TumjciB32c6/T3FkXCKFYCyE+Z13PKmGNPjc/Gstx2eyVuXvr0hmuJwdePO
CW7b4jVKJFa8AqTluzfOUCV/WTkHxA+uQcUJPRXySSq1XJDFu9z7AHdR5M4fNL72yfvL9NJgYJTz
rcytZvol49wxKgSKozGLdT9a7dnmRPHAxOX0eATWdSm+UMJ2gVTXSkQZJEVRuHgxv6lhWIbrwFvD
1bdgkB0DYnKqp5vfymv58fY0u82586yjhftxooakNUKTJZikc4jnhrAktimK4JBQgs4cs6eqDaBf
wrMOI8w/0Cq8GEIjqWxYPtTHs8Tte8e517haGUjlcKALXqlnNhRbOHBTUItNRt+tGYRUz8fu6VTs
SXHDq6MzvJXcMLFflHNc6ecw4o1sjR+ecl15GRlE2KHxVA/F3UUTiFPtk7MHEL8Q66WEOQDxLy/c
xiUq0sarKVavoho3CUEUHTRWy3rr8HSobhoJ8pjcIAiQz5Rg1nWHOAsYxgGHr8wTJuBrqHRTLZdJ
LUyOiBfFfbts793dLNTKg6cotTuiDlXV2yPkuN4G6lV9lOofqQlMqnK7zO0jMeIiJRPQYsWCNBV0
aaLwKJm+CjwbfSYxsKCCyoGawjU06Dp5OlSWExK5YrD3dNQksIcsoDtX/Sxwu5dmT1Hc6p129MY3
omRfKkWrkhzfiQ4i19aVstFYqREVn7jhayo6DtZBHsMbmpVmZrvIrwTNn65oglditrpzpycj3IR4
8lUpdfmEGsPS7wYPERS/FbC7oS+KvJUv+dPWm9lnFgclp5xWgVKvCxuLohrNEGJscjUZMO8nos1n
a6V8uM7OPe7KYyuoYTki7FZJyYRsWYAv7j2kW6/Kjdv27ceAnJHSkpuNxch/Uq7D9VkYIDzkU7Eh
zc9ptkctt5MvtMPDqaVnzq0kFOJgyXDxye420FTeJWSDop1RcAHM1oAK1o21ypGz93x5uN8NLAmv
tlSllVw+136s2v/ld6FawUS9gWvaylbRVdNvo4mip6NWcl6R3OL77IW61itJ8EtSlC6DdqbxStmc
BDSZtX7R8kWXYH4ZPg9RqGhmQixm0ogNClhxYZEVlFOMOPSmqxNSW/r3njEaJpHN1juerWhlcJsO
LKZ6nYpL4yJucjfiFQfPclwbxprsYFifOGfNaYrCCHm7Msytrg5ESQ8CgNKBLN3sQzufFg6LeTxT
1LHJzRYmbG8jBjUrv+REqnc+POr3yDdwmFr96n74zRVkDVkqOY+DMsgUK2HiEZmZ2DNrZpzg0EVe
0sqAhi2daJLSU2DgprBEPwxxDbyXxbQOzKQ9HDP5TpkcYz0BSejmZq+EMw4ivOhXXRhrtpoAhRKK
IS9xkCjB71337Fw4muEkPTioqcxaxDkq8uDyPs6MLjD1XHU1PrDQ4xCQS0iTE7G5rjZM5WICtssq
l1yJHbO5IIFkhrZutb87/QBW9+INVUZo7jBLPtEKhFyT7LmfBllHG1O46t5Oz+yW0ks+jsRzvtmg
ECPtXTmjJSCEdopzFrVftdVEl0GBZ7fAqrMYUr8VtsMDBnfdVrk8A5M/d9fkpHUeY7R4+/SZoZbD
bqSfelGorYne7dR79SI3G68AtlzYHjJ7AC7XCESughWSY/y/1b+wR0lmwm1IQgsQw+dBaCmQCv3O
9ZTu1UNMZuT4W7dS6bMuGQCNyPXJnFtp9X9fJsOqFtWKM8Kdteb/1rePQOeixlME/bCn4cq8EMJx
lkEB6iVzdIlNbEQiLCwCzbfILu50AhMPGIBDEVS6X3Ji3b0eQEKrPocmLuvg5ieRnhbDVqnfYxjq
fL+OEis53oplEE/IBSjO3L8zCj4rFEeCkohw/eLgYC4lDTZaSG6LD7u4BIdRm2G7IkWNoeECm8YZ
3tcqm0VIewMUkAO9QCmoYj0NRI1PEUoXCmxTgvEXhR/jogyWgWXiuCrOfHKpnV9Lb0YKnmZGeig0
lZWt8ykq2ci9n92Q6iHozMKCD6Zhou6e6reMb4O2aUhc5JaWgh3OItbaHs0PY3eSRVSL2zR2/dgk
AJYxl3S8YnXj0lau2FmQJdZPqKC5qctbixt/6eg6/gHlQ161hM/Uun9YQgZQpAXVf6wdLNDzjorO
1vgg5cdB9JsX1YD1VlbHiM7OoUBCLHzAz7cCd3e4iQkdoLbu68EZt0pRcrMZZMZ1R3fe5qiyBBJj
4iDHAKgqQSYgTufblt59l4sAx6t4KQdJ+BLdBwhnCFIIKnFnPmkkCfHI0swbey3w7Ic88Hq0ye7+
ODh4fzdCDAAPpCicw9adoyeuw7LlbVW5Ce7S3MeicJCaRjVRz4dI0xuFuNlsSukmJbbPyvI/1FoS
2ckacX9cXfP6KnNaZ7jYeF0GcALUi1JUl6rsD80keC5SzDTbX92U45Rod5Z6qurlrAR3o0G+H+XE
JN+OrbB4XFNaVYam9nzYCC1pAd+96l+/2EOrCH5UpptX4YIeHzVIHF22Ll95+1Fp9C1UwR6jgPIx
pYqirUBlDSeeaHHWxvyn3HdQY4pKWQG02cpQBx46sNdSRwBOoMUzxE1g+j2vAjEaipXyMumSVAuA
l2iOQ4F2BOxt9bM7hV1FZH3LosDdPnnpH0DODTljiR+wRJs1HUsU/UF2O14ccx8VzegKibUEu0KJ
phIn6S6S/ELGHF7BAaWBRzl974NcxZlz0ZlttNh8kDCUIql95hSmqwRiWvXyI6vS2l3/X3rZ6C0t
hptwCfbBGnls+7GU81RrpWKx8jSsb02oTEIYvtoax/6zqtTeJTDLQHNc1pO67qcPOfQCUyi1z5SQ
ER23YgOsTg5dC+ivluiAE+m1MdJSQvRsnzJQ4UOicv+PrCuo3GIV3+46TMN+t0FYsmCVzUlBv3LG
As8Hdvudz0JTXNRPXD39PpDe+0eDGgqyg13KWyn7xyZWkIPYQ2ELWXTBlxYt82aGBcqiF9wFiOU0
ZR58ntw15mmWv3hUEcgBtbn6rCWY3fkTAMJ7WMXOkc7dBMcftK3tCZq/Xjaa8KkM1NBgpgS/9Gpr
8etWOQsrlGEqsg/ogWwnALsJDqYfVcWITApEuIQwVlrBy1SRXpfxWdFLH1OD2Me40yTSi3JRJ5z9
bfgxcmsWqIsFXHpkv0onVvDlsYlkt5QSucVU4KDNxXmDr8wZx85yLfttuqLzjAm+lqw8d+LtA9h7
qnryghzYiCaj+lULsJh3bVoddRLo7QHCmx5JRKfS/uoFccZCF0HU6eejCaRY+CG1e6cTxtvQD7kY
OnZd9+2gcypG6VYa43EefmUlonI/aDFJxlKi44gdpC7+owzRyWuU/Za5oGSC1nPLGLxTUdzr/EKh
XXavp0OZy1s0Tln4yGIK3YJUMh0DraxCGDeb7p6F05M0pB/jXXHvbnqGOMpcmSNnpGjbJ2Bhcndy
UL33zWv41OSdbHNnjisa4hsUfgBrj3uyuHxC9V1vlhJZfN7ML77y5Qb+hABQWOgjwTHHu0dl0p4r
oYA5P8t1WjfAkQQl/gJWzUDm6e2D/84eneEYoM1wk9vUuFB4qUK86jJSBZ60w+xr2UFYGCKSnvRu
wxk2bF7gAr7+mjCqYipwofGd4pqOnRd2r8mSHi62mClNMUClI0czQpBvgnC18AMk/KzGYoaMB7Va
BYdALAv7qCZNtkqUBJfG/PO519aa1ZDVzP0qMBoEpDKoGcg2Gef7lVwwuaP6PI5bUnLg2sYxgvzn
rxzYZOU+OgaiB9dOrjej/ShHAirPKljg3VLQ0gFqqw0ax/lvcL/LC63mxwee4D9j4Q9CsscrnNLU
HCjQ55i3nuHEhlqGLShzjgeBInhVxQEk0fWfQrWH41cZziJg6+ViNwfJpV5ZKVmGyzyBms2ciGhy
gfjjlTY/rvUk0UDOchUO3onDf3+mypwgq0VSgoYNcSqZDy9PxY/hUeHnOPciL+bUV2shpPTs7RM3
951OHqpe2Wwx12153JzbIex+XFO4Cj9JQedu4X7r9JIX9p7vD0dKG5kd5Kfltm3JUAqH7ezuEDvU
VQLW5wI/aHiQS0DaECFmRAmK1LdUAyt8hZbjgBLbwYGHYFndDFfVT4ytKAx9Bgo8qaPJA+O88nL+
mCUSMa8M05q0aKTkDcAgWYgnr8cmaQGti2Y4KpFTGUCpTBrNujh48nhK5fVjq6zkBARdlHmqIEyj
N6TaIBkar9FKQuf/jTyulABKUuz4c7TRHRRy6PGRdkMCmjtMGelqD8Sjgya0bVmXlsQsUPmGxXbI
yqMgmaLbCeN3SvSR1JAw33YtPUUcBAFfZyBEftTvsFRTw7eLzf57ueKivckJtfRxDGBh1xrnpqoE
bjrur8LOY822B6WikTibvo9hmJH8kTXJYLKgj2cduarsNffTwS6pk/xVW5qW8u1IQn0W2x5re1F+
RQBeW9YJZrCrmf1XdqJHHnBWmVF7wgukL6XmWAyep4GANNyBiOgRTwEqGNG+BIZi2k4rN2HOpryY
W0BUyZp8wBNmMvNGr3hveXWelpsN+/GIbkfEozdTUjo5sR9KhC/jMYF0VeQsO4yfdU+WWeOYb6ly
Gr8Piu+9SHsd3db5boR1NVWYpU0A2ougWsGt60pypopOKi98YHdoQ+2ueExB3YnuBME90tJGoOF6
UZ+IR9nUjZmkzoe7Ja2+Tx0ivSf6/LKRBcerNw0W0CMJUNZjUM1j6kp/Fyms08L3kPdejTH6tr6d
cJGF2ZD6c7RwmaCQc6IfS3Rr4ycBXAdk+nnXWUQfo/bRydN0sNMBOv11cvPV8HkJSNQmHXQX9nrs
JH1A8pAgLPa1lylMeRYLpS9TqI3rfrOeNV7p+ujcM26n8n0yo8A4xm9xHHPNbQqGGjWYkqqU8+gZ
ik8rfl+ea3+4DKxn1uqxk5QvFN1j7g2WKKjJtg2iVGHW8UY1Kr9pN89ysKt3K0nQs/bSprPS50ti
8qnJEt6T8MpAIiJ+fbTZy6fB+3vZLFfDj+GLdUNDfVRox+nggyr0M21YIeHbGZNwN5kCD0jW/+J/
eJqewNolon97VmSBkKwK41i2UBVcowRro907nrmbSEi2BOwEPYqyhihGsh9Q68vaDKnI0lYCnmcB
fqoeOY2Nt4VwvKH7midZEF3imUau63jM9NVHS5QYxbBxJVwy0yXYzk7MZsBwPzEhbkBSeeSEKVf0
4xmUBwV8HxNmiyKKca/8VrNSDdNEUV4UzJfhaNiGIQui6CLXCnsESjHDxyM3HjKz4SuYxzaVGEzG
B59+j4x+GqCi8nByVXihVciwUfk5MIUafqIF+6MwISr4wLXEFU52C6fAepeHBAKklAKEd7QAxEla
EzEc0J2vqKojiPVVtnhG2JsnKbB0tD+v+uuaBaeyVH4Cak6ZzcQgK8HhK3Mre/Doa5BgeNR7Wj1M
Vc5jboWTSaMS0Jtat/xYOGDk8a1rDucisn0w3eZIe9xm4V/bU8gG5+kDJyGwW3ztw9y7AA7rxNB1
8SBn1T7FvKFV9EQDe517Mqem63W6hgW7EhV4w7PKGzQaBjydM2TXwgSblxaUY4S0cP6CQcvEZmhg
HUxgMZV0AkLqZQQTgAMo7rtwt8FXggVCL7r3Zu8to5Ud1Hv+BKoMA9rvP1zZFfcfluQZayCXWtvi
9BFjaYTUDTCmlahMCLhWhiNORzip+VsW7YlvViaSPyA1qsvAbSz8oYXixuLsr7KNJXBgxINvFXWe
mWC6JF3UzyRXmoCdRWIcXksJRHtHl4xILYxTn3EIKEulmC7sGF5GDFjkLB1orLpiTsDd5TG8ogV9
X2UzPzLtfLPbS2haFDr4hn4Mc8bGC7h4r/xqIbz+a/bPngPl+Edkaz2+6ZgFlVwe4MZ9P6zokRta
qLh0Lckyg4RO7gk0PfVaBp0vg1pCEPvW10iHbMS143MCjCXjOWeaWH2ekedrKiHtTgP6wzzUMN+6
6vozt4ikFZIzGv+XNIQaZXhhe78L5xGj5/iNVWAqbCzBrE10SHZV0eTAHCMhT6dvUwgc6nKbXocH
erJjFHcXpkkZFz/EmTpPUxz5Y1SPKEoccIKs1kCVZ0XVBY1k2z2AIyDiwpayQ/byxHC0Weedg4GS
ac4e/jtG1iPr0IxZEA5ydTlxMv09i6Bqd0cl0430fSyrxavaPPjsXz9cHXcCmWTh07DVx0fAoSXN
sLz9CwGeNGysZpMrakDzP//Cj86Bm8QSd3fKCfOF8EdPjNlCKrosw5zKDCGQlzWBGIJfCHOUEzAb
4ZcaP4gPfl5PCyAzIY1/ql7O2L1qj66QJbyfDhNQXjueI+ldnSsqVcDA8eF7UuG7PK5fQKLgy5f8
zU7/d1MlBGatFQWIzanytUZxqTFzweSHL2jJ1Uy/SCWD4w/3KolU0TKg01H7tBf2tQNt7EB38fEQ
c3Tlpd6Qo2J5rFBk8nCHHLuG8xxcdLzB4xOhcWyPWwCpc8AIOFEYy8MeO3hzvULGSKV6XZG3EiuM
vYu8O5R4Nxfv0Piga1EPkOiFvLLWSWnvxjUAOPo18xmAsciTAhVzPpliAkKNPjTgeHFtSRnaHYi1
aIIY3SazkVnmETiKrddp0gZnAM2cCO8Z6vNvakSG5fRGTXAQkSFYbVQf7vzvEJfFi6OHfCEZiXhi
yW+B0f1cHJkSdcrxTxM1j9TU8IqBQvldqhrQpOEeOkUuQFFPOsWdSJMBlnxD7KZiXj3O8RSnDdmC
4vUfucRunkEajyH6V1MQvKIQND9d7xEofH8g542BfRT8Sq8rh69oxAXWkVPy7Jzs7ezfpqQDPQ/t
KtPp6hlpsp588PYShb45vTmdt0BZQyNWwCZ462nxIpyoNp/P/pJFPJom1CieDL+5bpkNhBSss5X4
QcrGNvBJ5zj7bfZOMkvjhqNezdvPX2upiScKt7HGO9fzQ6bXEp2BSibqoTm0JMZ4f+J25DAQMA6u
I01OcKnYLkfzX8DzMotI6WlK48eq2UQyd7NQXj4CuTg6xkN44b6piqFsTWCp1jCbHFokcEhJZ3R0
sAKsdrRetowIfUGoZp/4lVdMg8VTk3C1wgIIVJSaVTCinyVHOBKlh9OSqrKzha/fgIZafmI8W/z9
ag7cT5e6Qnw2SV+ZLmTHw5XALbhHiSCXgVZ2xguN82cB+dBcM5ALQcFBsbJYw0IIgoY7r1cyejwC
7bC/8sH1tpkUOFlVrmHtguPMr33xO2jFgRFny/Mo5T4FVFVQRzl1z/lprNYzHUgPkhXKkS4FibvB
XLZnB9G/odCPedSffvRJ13tymIjGeqGyA8HbrxcXBlmNOaitVb5+3xbdhABa9754fuH0nsbGRgrq
/czupH6CKGcHNPbWLiPRMWq1st5HwMZcJGSVl70xvaIg3O/pTYe1XYTMwju451thh5taLygvfMGy
hhXDFFN6r0RkkKZHDNS0inETBjVZCPFNKZmTRcn+5M+24tHKr7qx77ExTd0wa4bYPZqzQmvkyjPL
B8Lgpevue4j7UgyjhZ+qbHwusXxlRSDAp5D+23Grxr+K6vIgVILYYbRmPuhWe+do9+dxEgyYVZE/
5aa1+61SjdzN/Q8g0po6OU2YbI4/F40i0vM39SeTgsjLYSw+198PxFR8MvISEmupIVLmDflVce4S
bUSuTnRWrlSIX9wvC0upNRu8VZyqCZe2D+1K/ZIWA2CZ532RxReX0ASSNDaV+KCrAZcWts4enoiY
GQkAIXlvp21MIdnD0/WmYb/jEdfuQw0/0v2hZgC7U2XJaU2QafNni8HXbIjtFOUwdHsRHE++d0Cx
/g/khwILU0Tau2ISisVQDZz665BAM+/YoTDnZ6NZRttBA1uQW/Ye/sDCvJp4mbXiE4P7Wc2R4WFt
ZnFjbKh0Ov1OY8a/mIH0Y0ioxfCuiS/U/wRPETNND1tNUn0Rtszoe9POjaJK4L/m0Zjp6Z+Ja8mo
KgWCeT/XVlwynx6xGfpcOu8t2JaFJj2V6mEBlqV4vPj+gBoeXEm8kwsJLPg9lC5duk39KqN5gI3s
ZlT85DCLBMVx2qXDTErMJPmySLVnbeHoCDxUYpAMvxEPiuBNdUxsggdltMyHDwWsCCIpghoyRoGV
31Q9f4TEp5ouLqOQcCtsqx54mzBFCX9UrM96N/rh9748lghXhxjrPUuMTw4Pvcf8HgdfFouZBmdK
a8xOtjM1IQvt3Q3eVX7IEHLrhASQVPDxAEmZqiPrQ+wtNkOm3BgMYp7zk3nmt8VT2FPnxHhpgxf/
nT+42hyaDKq0LTU/Gau7u8EgVmjTYPzp8+kW96H5prMeHzzEPejEKn52RSULsZqe/MFvhub6o8NK
/zzea417exwQ2/+WPCtXJWxIUaaB0Kx05H+vN7Ygbr2WQXNyLg+ou1UxvAJWofr+LBlRBBdNmKA0
gt+/Vef+3dTDPp5aORBN7IcZpXhsa3yjDZGgLDLVVJK1sZBAeGjNQsYv4SbSSnHrUO4L9ItNcUd2
aiu5cUP36bdMFTiraIP481gzanxg3JyiMJtJJiY6HEAs1jTUh02n4k9koNgC0idW5QmS9qK9/5wn
4mtGr5kj8ZIxnQnAEGB0ehqVjTK+g4qrzaXrSQ/4OczejSZ80fKt+IW5jmwlJu+MzDIVjnZbA0HP
rqzOFRz6XKnaW9iO+6hXgFfyq1NI/qO8pdMgKZplnIHACQjqopbGmUcMK3PrjlfEiQV55DjyS5Ro
SSefospbEmSoSERcwTrBwCW9OAXhFGn6hm6/PURgaiaz/Xtyfwyrx5wvwQkP6/T9M9KdIFA/TIjW
jnx7oeJdgY0tkXMPT4y/Rrx2yG7WAlUJjf0u9cdAudI51DnLTCIa2IzoPjvVLTM2htny2XnRnnNd
d+4OJ48+DXTZAux1CGpKOjsru2Up0coM0/KWqgcr7fXK5vVTX6pykAbBra3E6/PTgebcgEESrf51
lHyRhyb1l2H9yHTKs0uEFRiIe3R2BTcyGnsnXj9bQllK+co8rUR4J55PLtMRTKanBzm82A6FY1Xe
PEk6ak3vsixrMWiKBksuSNi9bb9lN45KCdRNjZYeRouaIunYD93iTNBcf+DbVLtTM3eZkj9A1mx+
WvyxgxPvDnmjLzPYXQxsYmKX3jVHy4iXseQ7aPH8rZ5vIg1KUFzWaPOelZtnlQg+3nUHYUqNWBcW
CuwTc5gD/PPvzuI2Vaj+Nt0aW3fWfNkrDW+69pGEoHGzg64x/Z6VXUaeo+moYS4BJtAEKgaCOTZF
IWdygmSz831xviAFcbaBYKeh+aHXpzVwtg3GzmUjfnq/HniirppJhCTVaulxRh4jTW9rAyphlKE/
2ESBbgz2TBIEzrzDTMPSunkhIlJD7p3mWZmfGV/usXcp7AVjUSVA6SQos6Aetk33rNaOHbKWg2IN
5WbfTc6SzjgHXirxENdkH5w4mzy8m3+Q7Wxjap8PQFnjreaUAg4+XaVCbctLfmwhewF7US6o5x4E
nwahk1lt2RhUBgg3cb6MKKp7i+3HcJbidam6UsOZFr1R6rucLy7V0oV4nU+fnm2/EoOHwQp6UIlo
m/0jtznBLfwCwIDwy5YyQG/FcxFvA7gO7OxHLp2u/nLKnECzIFPgKeOU2tPwHqpv7hqVpmKQ+c/d
fOMeODxOG1+jHDSyrnnsaTXPH/XyQDwJw56RWdPsCXYKkKQ5lmjiShd75pvSAMhfeI4Q6FNFAQMV
a2HAu3TZagAsLtZp+pfvDvDp+2U6x1j0pyvraNCrDrbtXVUwbrfMNugnxdd4lSKrR7MfFwZAEQOP
PXPMkT+Wj6OZ4uvaHtsWTolB/9PuuobdoL+wDNUmSNgEPiDURSvuFOakS93/GpB7iHczg1uUE474
0k1kybDiJkFgmiQLRkG8CmUkIe0Rd38eJGP94jfRLlgMrUN8bftJd6pLh/+w6L3qccMjQPyPaowY
5zfCJP3Ez0hZmL2er+ghwwvuDcq6XnO820TEOtIrbjfRgOhnb/h1AmyCecImfqV9VfkMFJDEfaaM
uZ881k3EpT63ViaoSjWroefiyJztv9/hnW6rwAC0Ok8lAAZO9khDo7kFU/eXFOVOLZrZQm9rrURo
Kg+2Cp+vmtbGBm5rycsVHxsfJ9POqVaKwpZgZEQSE+Cp5utdoWyFCCI9ndRI3hDv2LGgkPsOEfPf
TSTvgILTKiREAVDgV3XYy5uyfBYVZODSsMGDfVAVforddFgpQwdFLf2m6UnBwk6Tj1N08JD9Gtzg
8Er974rU8RFws83BqWdDa2msytwuR/p3cPgVn0Glsv2IbIqvpcFDwJJZ4dzUB2Phh1hyKR4I/Aud
mzaHjZr0ihGMnOz61diO1VuDDUw6EgZNVePxzTh+Tk+3wP/zo7ceWZNH0nSM8fp8HWORWI4R6lNE
XV6ns5C3fe/9eZqo1VsjH6Ke0xZOiCSKSoLsPhmcPGWtQsLInUuJ5pzaHPjHXnUbpNVcZxAx7VDC
e3yytisCbWyj+9d3SRmtC7ebXGHA2QjsWHa7HqZYV1oDzOa3GcgT/s8lbZ5kv0zSlgGUZ64vFU/i
RAlOcvbNuvFaaQ9P3zea9u5wXTga+Hy7mHUvLQDYU0fiG/3peADgL5Ze21nEOYuEnI2RQUZ9pcBV
bQ3L17mWLkQRi51VOc358tvWJSJsV7ZjOdjDb76JOMr5KNmUibalgd9D23dh0GUb7e3ciUWFkT7w
EemnCnniRtJ5F7khJoekg5k/cH9Se9Nih9x5Pl3Sgk2BC6/7+X4xMikM4dtpocAo+2hxQfiHQbw9
oKMbZBCgc/rNkhckQZjYkA2Rma1dol3+0LHWGXGtvRfnFtDJ/+PR8MAI9xOwnQlYGcvCM9OGllUK
UFMBcR117XAhD6hAwVL8l1G9qDQIpZYIqfXN378yd5Swe2pZq+ULuGP5t60Jb4H9seUAfj112ZX4
5ePQgbsH8zEqYmA5WFKDY6m61FjMt6xnTKajR2FZZRH6BKcLax1NFNuZEas/NIehxJCrlF9yozXA
1XDsxncI+y5LQxvAX5/lirPsZFvJaeAOV0bEFTnS4W4ZpsYq03Xc3Lxbc8OpU9QEqjmqfVazfq67
W0siMLw7KWUgYzfocEFLBukPRSsQLEguZQtR5Egv6/qgiNyrxr6sGBLZxUMrO7Azr6aAN6YsrAzz
tf/N+BKXycA4X2Y9bt6yO7RP02h4oJUkmzvKHy0eLW0TYwI5jV3m9CphF01teCEm0rBI7BfMWJ1t
f345Mh4DsppIN7t5WllrZn42T3BE0GhzgeiGj5cftlS7T7XwCfYO4iJItf53sQRVmQthRoSdcZ6i
G3lo0PhBCtasBfWYX4VnncdpbNDXsIrZUlY4wof1maQcBO4H2wXnOadhmCzsB8WPwnFGGESbQNG2
7MiMzsKPKpaQE76Zac88+GrIev8JZERHilJyf+ANQ6ZlwFtTPfroW8uYvLc12r7JwilmlqxPdk00
F5zB+Leos6YUNUQaZVbi7EkibjHuDMqFNFAdFCsxatTN2wRGSSLwUChWD3PNC8xaPQhdFL3MZgWy
CcNoo2DOjw+ib3PZ+w9N+dTE7N33CWRk2CkmXqzEjze4mRNaFZlw1y9evY2lmCk55S85aM14LBQf
yYdRw1IST9gqax+gy7o7TGlqIb8oR3SPKk70KL6JWuVYCGomodeklvWuCby09BZfjA2fhU6rz7+l
qjAIMKPa4UGqlUd1GE1L00dOmFJJ4LCfXP+8JbJZ8wh+ip5i+/eWXQZ5Ij7GQNgwm3IK1MU3iRCW
wdpb01Kr20RQeK+iiujJzuuuU+4UdwIPmSmO3RbBmsQMLcF2ZJqgCRWhvhGgkm8ByGLbhijbCxKj
PCprhEKqdXTICiwgRh+ZCTDGOIQhyeLIBihC0BhQIa8CWFI1FmXor7BoYooa9bARcmj8NS1L8LdL
MNm6brSumXGDc0KxJNZB5WEyaslgJ5B2DDbYoGeCf/LRRfFmQu5ctMj3BrAqXoQ6oLU7uZlXGSdt
6jzjN5SY0sWiKInUSyU/iji2/IzGRPa4xACnlsg9TsUZY9BraLlEdxil8E69elx2QH1TQz2mV4v8
7D8PNXQPMbzlOiN5deHz5v1bk6uBjXhXV/fuakDwyFIxRa69mX+mYZ3HPRoG3LPf8ABRizg4e1eV
jYCyAw0tPQMbCZ9GfxdV6qGYQDuF7W92bk1+kSZ0KVsLi0Rw/nmFWYz7IzmrhhYCVRRE0EnSdlqh
wsZNAtFMdOcx8pUm6G0q7/4n96UHC1lb/oU8fIL0fNQO2TGoYaC7vhlCBKsOin+d72DJPXGF8LE6
pts02XBtdRfICVKfyfh7vf6VQHXnrLE0oYU4n/FqdO16YHSrd/brvwi0kW0fEQczfmZnCbGwrj4w
7VVFTOimlvmp6eU4rvL2fwllGx7w4TzRQzd1xQ1CQz+oi1RPGhx84rC5cED9PvwPiRTYw1Ma4qwS
/pDLdS5l2Avlv37kaeVupGtQ01XgmauqyCRgM1hDJzFZ4lZwec93bFbQCBxpgjBjEcFMyt14x3HA
l0aG3dhX7JEsBzsVt55luBhNZqFwGKvUbU2PQm/CUOKTcHr00NAmQUyo8D3hq+R7PLY5fVn0xS8E
duLyaf9n5dKdFqzLxbhI2XqVL3gzkh+tXAj+SLB8appmZRnPCJ3l8cWyHXA5E3n897YikKFgJjgP
HxIGTBMMBoLnCoqM+OXnpT9n04dMbBlVO2eRVtCB7CngFGAhFVsIvtnfDSPv2aZRxQl4jRCdM1oF
OFco5/kmQ1p/ynVLQ4xdkk0P/bKPXMtEVRpIAehQhPNSv9pc9kyiGvn7G6zuynZWt57MXt/X9w6m
yi9cQz2NS6rxZ869aF4XFZE21pb/HRoKgTRqAFtrJBLcPOi5bx/ZQwr0MVVETZH285rfiAtNMksL
O3Rcv5jiFPpdGygxVhZQNTi95PWX1J5i2w+CNTK3jNhKCHUdzOcNLH16G9MZ1IEmOKTwWrUMQvVA
Tnc2q9YSc4vggQDsnMV/5sDV91TAy+xT+5O7QNWZ1pv4P0n9mSataYQ1WzWLu12UaQCSy/NvdMYi
SrgwCTrBEG7RZh+D4it9ll1vInShH8IgjC6aCdBYdhT/TqSNB3KFguiMZobsXTmgY9aImsrHrdKX
/U6t9GJ8GFa74kE4RiHds80cUAJZ2othvcMpQ489nJgHxFa410G5668NpQxAxE0S4UkkiM7lAeN7
6WBABR3Kdbo/qat2Q07VT5PHSBvXTko3DlAHvkGnY9+dE1GnqAqeRd0d6GWEmBOKQaaF71F41mjz
R/ElTD8sykvuSNZPd92/L7pzB4RqoJQXe7tJig/rqhVfw8e18oZNTplzo60A+JX5/ttxr0WRIvC/
GOcg8B1R7Ze3zK4iiERcG9fogPxletd+82LQpOzdJq6ZbNb2HCV8DPPUXEA4X74pZM/NduN32uqG
QRspeenrTQm4gu7qNTOsVbbW2xJgDwXKc7XrqUGY3ybrxSo1szehtkSzmP7+ArJLT0MWvId/V6d8
Zu+5/G/hC+euGOEDpHd2y+Sc0Etk1SUBNkvX8kwPGbhp74RzGI1xeqSGmizdTXIM1PMcnPYu/joj
AmM6BzTRaQLdojtnivEZe7a8S33ZrtThHsVTMoaYgAIdCen/BA6NjMJ7HOh6Xtj85FywObKxz0NM
KhVomt8yrrMkFOga7hqNwU59tsILJwg44K1iCy6vilS82HfQhSpPknFtGeuOOZO9SgwKgCk9x/Bb
GQVTIdtCYmzgrBKV3LH/N/cVWhClmY2LquZl2AskbE5zKczcrP1psm8hLB86QXhyMoxjAN0zkL4P
l+hEY7DqTL05TzoC1fvyx5xZf2x/7xaGoke7DvyDXHm/kmRon5xpibVikbUNQ1sQWM//2djIrn7T
O5PflyN5JhiHDK6ibEF+gQ7I187hFtHmrvlG/daCaqGtRKxhbEb1cKBK6Donzcsp42THQwppGpHo
fSoEQWv/HjYbALaFzY4nbcupv8syTbiaeM2B1bpdd9Za+Guikltu6BKPYtigWTMhheMAcNTsRYMR
p7vjeD27Et7ZFI+E2CLZyFRKVx/Sq0QuwnpI8V4mfYNgZOh+6AYqdp28XRWiCgyW3ZeTu/yCzGMd
PPBNWORNQXPFaumE+3OjIaX/2SDzT5J8h1XYEcOBINB5A/NAS1rPq0XK2/8mKh6MuWDlmocNzf5d
GSvhgaHykrmCcGfcRWuvndN7iXdlJVlcZWxS44cpuSfFLr2ekjkPtzbMwWm8/0wvzvJA+IpJBv3K
XPKT40kpcYATUJPgI4GTWwHNNcDnwpZpwyhEobQk1+fof4gW45jl5yGEhWOGiKSxqaZ3KwGgvxXj
LTMTgI6YDGWkynVym9EZPute11FfEfwGFuzY9yc6ITB7/wZf0RPdWUEwkfVTOOA9fBawm9i1/0+Y
SPU2jDJH43HjCxYPzdR+8zxs3FXn7+Y1OIHJi6FFtJRiIRctw1AF9d7mTBcZZJIUsRWSfNcSO2z6
yERwimSj19Bz40sN7I/LePZ0SecnmnXid9iazJJIVs0yrsPp0lyvvYCW47uNaUyDVWAhUI50qQXc
bpijbmPWEjQUPzFvs4Ab+OtjuCXWMhbonjCvufoMBqMylF9zrkoMX432FGISIRtCT0fvt+6HEEQu
/6bBrOPBJ6Pg6xQAnAyZodvzv+gyemu9bedpsz/dJripXCrMITJSiigedn0Nk8ZVDpiH2agsg5n2
86mQ9Th47MVZ2pg6oEZvH0Ow3L+blm3/7Q6699WrPRXhWJtxM2u/+twbJDNXfcU2Wify/hYxr7Gj
d9exlA47lMSqZyXlTvRObrXw0FxZbn9/v4wWJfMpmOGjTifZsqgy0tXNHbIQI+IW6ooJF/S6cRSk
QrA9tw+9MdboMHI5rO7Ea3/mm+I+HsN0gWAEkY7O0wB8jJBjUNImO0qcuvBP2ft+De/54kXgje8z
me10Xz3KX4kg2E4W7ecLD/OgzmfGMHZVAvHmozGGGBA1IcAHLbJ40owXL3Dr8DGSPW7WbrwIp0iP
kacsgxuhfxfzXL9MTGHFA1wW9DGI5yfvw1yJNpgYPKRMoRkfzHoUQlEpKbooZB9ngYVI8TKEMqaF
Ll3356OUBoKeUy8beBBiOdBn405PkPme0Or7jvRy1DfFI7Jr0+widsJBQnmCPY4Aous2g0AX8AdU
CRCrXgLn/aRJwMqhYRce6rp0pLYw6e5WLqHWt69QQ/09bjoP3iTpeNf3w7dEqqbSIojDG+vo6B6u
M76B1HygOf3B/7lpG/0extp/fLEDd5BBvctKEiNAGGx4M9RG6x+0H5xQsbjSoSjL6wQyOEk89wct
V1hNYiSGu7sZNBWa9XfWcJWMGkA8MlP5IVwmKlaXEEXeSBW15xsnxRa2MkvJM9cdFp0kr/EBEgQ8
U2PpiBXlTWJyq65ZaeoRJKgWLwIdVebdS+sIKRcFSabRGm4LbP88WFiXGCNpbB57/fFoCvDE8YHy
Mv2TwKi5Bt00r5fAAV4cPanKDWmuuCGBr6ICz7wruqxa5Cx2BTZYLolnokmXhLUNRwhMqppE0r2o
LGoGkGIKZWaVrevvvmA3nE/eyyvttl8LuHnosd+7ai5iVtWk8yK0LCJFzdTgOXtYyisMit6y2kdF
Cab3njJiOT5CyYqFdRh64nf8ruFApfKqHBLwdDWlC5QN/Y8xeVtGFSYfbDPZevmHr/FSD3vfzSKs
CxwVUv7C4vst9nCr9DcUIPqv8HNO1JKBjJSbtd0Rvhb+c+HEaTqi96jXIJT5puQs3qR3WqXfMT4c
N+Pd+MV+LB+m68F5haeGLctsVMUbp/Qjz86SIHKgL5RBwpmjGgfyyWmJVJU1xAVNGg0F3Ot3kaUz
uWykoG2hYrZ0uuJVNHYxBh6Cdf4hY3/fI5EnEN3fachMb7afv7F4fiBgt8Jf6MHmI8yoUGVOMsjV
eOoOx+3LpF4Hy2PkANlmOio5vHpShi1OtTJYounpowGS+fd3nBlqmLtk+ovA+p3AFc5XWGpHdypY
Z3866Kz4G7dPXlVvDgiakJ97SoqEODQRdmcJIIII+/Dlzaa30xIkaCuXwlVo7nTjcV0Jx40dNsAA
y6ASRoM3/JeuhWR2Udki6rGO+LIvCWU+2DL9B77bKlU+FRDVIi6Xpzlnl3lAQ/QmLS+0MNnnpOAu
2N8FArBHm3dPI/+H8LhCrPw47yerpaStmm35UT8dvcOgqYA7hON23tVX6e7CDkxN4QqwTPk4LgUC
eR1KZIsiThnH8qKJRyicQkdJLQ+z2NwoEa0eJatqDEuOkPu2QMkB133VXu8kHk4iALanRaLdoZP2
fV+flsNphgmFaGjgfDCHIXCNWxwHuWo0oLPhjJg61GxAzliFbnPhCdTb+uk6tdvlX6mtht4aEbfw
RnulpzUp9aOQcRM441UoIh661E/T3eDpjm9j4BrgTSmkfK8HnO0HkL5+V6O0/qAl/r5ZHjl5/H8S
qcDjr2lXma3jNV2zzhuYw+E8lxq7sjLZTgIDz9Qtb+RL6wh2y4ZhoTxf/Y+ljKfRVaZEvpIoArG3
DqrsGxKKnqfmwolAY4IQqLjnvCKUO/+4v6Krddw1H94B1xpatveN6sAlghR4zyTbvPyI3GtINruM
QKJgHeQE9+9TmAxI4V/TwFf01fhYEWVWUAijw6qbFrJ43MvYc/cWOw0u1ijEs8n6F5/r2ihEtFF8
cobf9v0fBPm90TthtG9/f1ZnR7E490OFtIq6pbDsk4ZO0ShqwEib1cxEm41n/wkLQ0cjhLUH1+Iq
YC/TMdwd/y44umu/NvkfvOV6T68lvoKUkF3wRiXIAOGJW0TRTCjqO5gMe2f1sqkzF+PBqDjQQ+Cj
VtZ3EYwRHEsIJd+zV5NYBp9Lm3Wh+vd13/YS9wPuyRahTI543rdXjZ2fGTbwp6u1nIg+UeHai7ag
cfgpZfN2qqtOzjXzG4vHuvrColhxUwD53wr4dGbR1U1IQd43ZB2rt0vNzd/4wPLnOI5rCHfmUb4j
NKCp3etFtu1v872+ivOyRELZs2XvXVC+ufkX4HScO1GUYMd8lTH8vikA70vtniJYfYWOWfcU8eeB
sZW1glqLlgHT6JPdHjg99eeWnPOLkP13318exQROga6s9ATImDk75FN58wp2n6+4yCNHkhrqgx+u
o8OlMGADNWEB1De6Q9WdsmRlc6REnGQ52VXHncXgkZy81xTcotZEzcVNQ4OjAfO+LFCg0rzOZ0Ta
JC5555dOC84UkM0uF/mGn/yH3n4zUYIR/y0oEPlcqc/aeeOyzw7BCH/I89EJn76DBuemwkX7pPmY
0fIIp68weGsGnDvXckMPb7HFboRxR9m9rIIai09/pb5u4o2mwdRWNL5C39r/V47WCr3EwUA7+KFs
n/pqz1dPaS9PoPxq1zumYCVCh4wVHDsLDtE1teiNtX7smiYIIYPiRtEk6CRgtYFgKqO+124KkxMk
G4JJOQ3aZN6RVgr8YuUVDSsJqRb7/2iiPyBBfBk4Q7aTJhaV1n2f9KzoxA02785HTlD917nyQL6X
VIZ469opNx24COsi91/Ews8lxONwGKnr8h5hpU493p+OqD/oL2NtCOatedOKUabos30JCJa10snO
aX678Hs/fTl5RfbbFZ11C/SaeP5uJteUvcHfWQauc7JT2aKxVNbEAEE86b8uq+E0/JJkfwVUZPKe
930DoOgwR2Iou2yhDd1HPGuv09sVxq3Ep3wPVkHs1QImKOXhcg8+Qi46BearjzTunJc2D+lQ83Zt
V5lonc8btbyiHmvBD9RNScrWQX+YPVp3uCvzJ/w9dkVFWsYx+q7ouKqWviiWdasmG0ekfWfCD0oL
ldsSKbghY2y7cKysYY+AzpOULvZg1HWT4DEbvDhXjnUlmLouZAM6RqHB/60hKO0F5aFH3Pt1UeHB
vzAlkgE4iMofjhHw3gtWZJFgVDWncouljihyRFkmNGRykFPpWB8oAeA6q7AParm4vNAOgUeab92T
A1xqn9n6HD+eUynWA0nt8ntItEEaXJ06ybFsAXdbZoP13bKYWqp4FmQZ9MT0gUXQ7uqgDQDGjQxd
y60d/sXDzUyggevg2XZUkn6zXvB+2BFiNVA5KeseY9vYHrr2yqoADUvYhtNmVQ6jAf3YkXxAZS1l
Hhqh+cIq19sH9607Eb3o12dGWST97fPGkYWppqrE+mgym5HoTQ9Q4GQ66/101kYQtOsgeK7TlHNV
uqo6t3pFtj0TWtPMxtBm6zkKo/lHBKWCoCFyR6F61HyCO/UiEPZ8gAVbzH3zFk0ruP35DfPMRfSS
nHI+TC4jatEOLUukH6ez1NJaiEeYoPqHRk/JPd5z3hDffp44JhVfaTXkExd32IIRlcb8XvXN9gtI
dtx9WQF7M/HMHF9MjIB5i+My6bkfebGU/TVYYzt3JOQNpWSAMQTBL7T2NENYdRK2P3ATVlhdRJgU
OUq8ONs8yozRdfoBs8lhLOO0qI1wizE1rTeVYCkvtJME4q8HjC+MJtKDUgZcmXWobTaCJLE+zkEd
+/CMESz+cdy1aALz/LbTHnQDsAiJuGM7LDInpToBW1H0ChiCuLvqlWvyBLGxQWfcQKTfWCSTLHF8
UbgL+Nw6fhNAiRqK28WSkmobh8O7RJqrTbuTKj0SKAD5m7R5OCWT3oxQDKAglTdTe2kasrnnwIao
Q+U5NRLHp9SBNLdbLLy3H4gnVf+ACGpclcAYJdoaNg4O0LfvZ83sSneM31ITOkjlDwyxgbAON+NL
ygget4KpWReteSItSxuKysRjPpkGsK4brgK5l0LJ+l9CoMj7FEELHwxuBCAoZoK5kJiK5Ole2n4F
nkrHWSSrTs+o5Huqpszsh9vJ+6AvTkcGnEn9rgpO5+T5d25ZW7GzdeFHn3/0d2o+U1CQpBggKGUQ
Ts5yZntzfUylAWbMKX4HcvXN//VnKjmF1jMfLgdpSDUV7mVBbh0hG2ydLi63LfEQZQB+1NkCz852
kJcmXVagDpOqLzEUqHBY0GdQ2S5UQeqC7QIEVn0DzQ+5AoAHFi4Y4h/lGSEeEkUTl3JmtvFx2beK
Uuf4LgjsJIOe2QSDIDPbiMwK8Q4W5zXDny5TVle116PYPq4MTPFY/7d6tIvp/hbpNgAqYbNJKliE
PVsaanoo/iJH9w7+GRu/7sx8DT9j1DuO1tb2I/LCAeQ/KedIYmil4/FZy8o37GAgEBRBofUIfOhh
KUl4bWhCHnvfeDz8n1Xui3mhlblbxUcneyEtNrSObWzov2bzGcXNo50wxpSdwpiclbIfZnwsHO4C
ObGl8T2v/4dyDhZsZQRu/7u3RtMSpQyAK+XqViqqj4ZD77VhwPvn0iUK8T+sIirumV1EQqgPTVIp
PyI3KeYTVWW0V9gKt5OMV+FVwGZEJyA0Z8nLC46Z33e3BdVpriChv5mdKL0VfNdY3dH5+a+sKXkS
Qv4OwMzu2VrqHaqQsdomrb8bmzpXOMGEGcrJjHRD4RML0hz76i4jBH/HpBL9bmclLcPQvF5r6K6I
HbR9hJs3A7TvyBuLfBGlUXR/VRpdMCIqIMNMJDK/K0Ke6zEgk4nyK/b2bQdosP2C5+EdT9N1Z4u1
030gC1lWcX15aouA0iWw10S4/ZwFwLdkPwbvq2SzHYJYO1VsXC6L9ZStyDO5gFUgEZeNevpMTwfy
Bk4i8qJ8rNOn4I8PGeSxY5vrmB5BBRtbyh/zqGmWzBbZLjA/ayIuPOOjzxZnxnXP5NsIwHY3naKw
X0AC44yXQaUAhIqWK+ew/FyuNjq6WJ4EXREjFlbfnpZEcy/aObAgmG8UrGDkp60ewj/bAkqX6d9a
/2QwNAglHy7jULXqBYoDUqpmhDA6LgTTf5tEAk4Uu9z8V25VqVsdzYRugjl10ox0X5s2Ct5/0aaK
O2JWFbLGgrDLvBmBjVxzkv6AiQZ3afUT4GxtgaBbuFpTUX4HSq/bozrA8t9m+eao0rhq2k7dp8k8
+QC4zmeGJfqAg7KlFLezu7WOyElaP2zmtve+oMJ6WKLHckGh3pjcaZmAPmZBapxkk6R4o+gCE/dr
Hff8qmJIhSc4Fs0iXWGdJLAcoFa9wjq7MP73ifNeJ2XA2bCAzJU9HwfqFnX/jgfUGXgODMZpaJnp
/0c2FZOega/5WjHmW39zfaE3tDgROd/0OZ7yCMKB/1HdvTCeKJW3zUhPEhaFIuXAIHxIpgwlybe3
eORYY0RlYFt9l6hcPchag4PRRped0za3ypWrZTIB6Buws0MEe6FA7uTfj/eBNyVD8oeG83EAwrvR
g4AZrB/wkFBRgM0vBSJVdNk/rsmIuDMzCNgIe/l+hhlrjfKXiFR4rrW0OQLDj7z5oJUza+UcdmOS
dwDfc+gzf/xCaM3KC2JrjaE0iDN1ZdCK0B4Wq0+MnPUNntgFYkAO1nBSGp2dE7tHh+hK5zVfJNfN
m8hCii5xmyMNTeYN2EIK0mq22vd9fmXGaRXIuGN3mbQbnRwFOwvoXU/Byk3DBzO2idCyvvWOUut9
15Waq9zLMonczig597+uz9HFnTmxOj1ZG/7x4/24yowviuvsbFXlCVEW1RctFch3rl9Wr3d47v3r
W3t0UwRPJEpGTk7jg9rXZwiGQGjN6JAfRUyplStMwgQ8OhmS94BNZBXXLqihjy9/XFepLDyp6/4f
yfRQxu2zx3R851UZmOvAyfnqxWxlNYFaOBRWjGjlb9W6+JpsqjZJ/o/q0ijWmM8E/xzDp385TEB7
tgGg/EAXoPXoxd9MFBXrFCra08cnf0RoUVr9vpcJa0J5t3sBV9rq1BID8pZ8n/UWgR65H3XrMcsN
6e6eQ6fxOwn6eVILFIfi5Z7XU6Ww3S5hxNdmLTB/itk88EZnYavD2XQz4ZcHmTjz+vhjLSCqhW2f
KpFN2UL/f3vX4MHUJBheZfBWRUQ8fN0v3Gnv2q0E8Eo3fLhdXzNcLidvDg7M7hLxorFqRkh+VhJK
XsJecRxu7wRj4I/58hgiGwEIjzQhdOOpN2k+pl3HbKUciobtOrFINicYjsBmYmN3mZt0MZ/tKSAl
XaWn/zzlTBb+ExDmS+adMEqqIJJn0DGuk5lc2RMn1brcGhFcAA79QMDQHwRwCScqtvYdlRazkuvF
09ECVrlIKGpmCdy6HW5WIBTje+CrRu+nAEDn2BKGK7Kvat8gXX/A2YluXAl2CWSW/D6MBu/pKr1N
g+DBXqeqzL/H+UYWCdlOlFGc2lDqAhf4bquL+ZHXy5vVhOvTG7xvryWYE1AXyKhwIY30G6wP+yYn
Bw6I7gf2NKMrdrbnxeBk2Q/dc8UYiJ99LvDTUq786soPIbVmcWI0sC3GBOlxcFuMNnxUuOCQQoVE
T7sGv8yzwHovxL2nL7qU3FPZmprQBZZPDjdrQdfO3C5gRMxDBfqXwVmLq5BDftfSs9Hc9sJrnX67
jOZY03CCnrH68QWxbuMc3OnLcyM6NuKSmxerhq0sNmqqK623qfSRGJYXL7rIxKYpf0rPkdXUNo3b
lXWFwTxhNL31hUevzGOE/d9zwAYRV7M9Vbx2ZD9yvc+bJRFbdlTBA4aEbAivPKwCzcY0jyW8
`pragma protect end_protected
