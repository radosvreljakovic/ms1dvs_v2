// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr 25 05:42:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pVaDVhw1upzas9xqmfqdGui4/S4wMOkgCJbRpKYPkyztJ6GcQL/+EVhwKq3cmjJp
cv+PL0HCJ4E4aQapaK8u9S1RLTqWfYnO6zhDIudP8sJL+93IzHaLj43j/uXR3ZS1
CX7araTqBmWhxZ0SjfiVNSj3sJOkFu0COG1sPq1K8VA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12816)
UUm5OcqkaEeznvwNqAIqC/9xmedfSPR7ju8X/jUMQXB4dSRg6BAXSPJ+uQ5mMjpL
mbx+HZILqdJo1JGg94KzFdaPPOECq3bSwH96qjEbccIUYtii8sF098wrpJlfmMFt
pY61vIqS/5eCNMPwATNYC3voSxXWxRCDiIINgKdg1/TmY1QxdmwVhbMBvz5M5WPp
na8BZlgLu4ksFiQ2EZ1bvcKNFVe1ZevYlXyingaFP86fF8Pi/bWtCvzP+TfXMbSh
7rXsBpv43aGqEb3CWnRFikPg/7qskGxPA/eRdhV1tlrsMZVszpwc11Tdd9PsO++T
a3N6OyxnN2+j1Fob0f9G3/YWexbE2cgGo1SutkOFF/xg/hsKp75j6UXy7T58IpRp
qaPulG4DAWDjJfk5dK41y0Awvgrt80/Wh9q2aZiQV/Hu859tl4ThmNt2AyWx0RVR
bhIe6VTBbsQ+NCVwTHE3UILjSwL9kbY0/CR55taPWq0KvVkRYvRqP1iblQwTg1vN
4wLT7uno2kukp2hngi0o0Yj5np8uZEpREOnoSmP0a0DLK7NNGO3Zl9u1r4EW3qHu
NAEN/Vwj2eYS5fZY9AZakn7mHY1n2bZHcdFjVMTht3hG02sHbtlVMuQ0bWsUnikK
m0/KjLaxLc99CIYQvi7kcJfdow9EBC1Y5HYkGTA1k+rbNv5dVvY1AvI767QmdxZn
lkP48/fc67fbbVc2UV3S5RsfP80b4yO22ZWhvipnrIEGSkdkcnKq3eaaQiPgmXrq
htCEGn24wuDu5BR3/uxwpvCJyQCLX5xtOB+EKArfcnCV/uhWWRDR0+JWHJmexQ0d
VDiwzPuceNVTUxDOp7OphZsDw5MGyK9YPMsFCaD08+DwMhTwdE56dpAr8wh5mef0
iVA2oN4kwuj6zG7HUyusRfd2I6jLfkBCDZcjj9tXjnEJccU2tsRxM0wHdKKW2d2h
tQV559eA4doIfO0i51a5WSD2z9OxAE1pRYp1ho7HxP3P4ae0h+u3EHv5qoukwm/R
RfxwH5hudBTkzcGOoTzTKSgYcbCEklQA28AX6qcatEnEKD1f0U62OcW96fxfe6MW
F+NAiAo4+Sa7uvur89/lWB6TLMEzHd+eJ/fBlGqAqnw45XQiojP2yg8SQE/EnT+o
Tt0IwHtjbOKy28TQI45K91z0GWIdyRvwEurDMPmcZ+h2IJr9Vvh0kqLchRJwXZqi
kLdGBj6i6NFMQd3ACI7RLWA1Zk7ILugLNXsHMSEcNxRp0bWWQZEDywl6iktf7A0x
MnxkAoht5lHuuGpk1pDL27D2lshi/14V8fczPF2fb48RZP3SwhaYUOOGec0Hm7wd
qUOcnLxnEmeJcXLZ/ZoEH3Alfyxn7UUBXpvXZOIE4p62db/yPgxvNJJSlAUwAIeM
hJXMeamvg5NQESucvYm6oiXhJ3xyxm/BZD7vU2hwyjGtzccgVr6y+mixSdf8/FiH
5hlt7ULW55HSOsr+BrZYJvi9TpZ0iI4zRMohTT9DiFd5LWVDuHApNz1QZUOVbFp2
CzPe14BrwfVxh6hcOp8dYh6kKMFn/AKJvkg2/HRDRSpt4Z/IlfnJ44pcwo5pqCM/
KKpVyv5Mue5PRLGf42bdqBArdeZZVsWDkOPA7wOFQqXZe9MV5o41hqg0ZUWkTYOA
XF6iVb3GCmVgj3sK6DHelGHZDeG6iPtDNdGSRodtu8RUHcjdnNPB16BM8b7SQivh
aZPRpeM3sIFkGLnjDTrHYsaukYY7E+7syt5dkFqgvVb3ui17Da7gxjTrCe8aFoeZ
d+s7MPRQVlEyO4NVW0okdqLOrSkNy9QSaT1lBfah82kpqP1vPwxOqlM3irnYHINg
v7zzOWxhGU/wy+VA2t2nsxEnzlXWpFj3j5PTGpEkbHnEQM1dA5ZvqiXHV9lTRGY0
/7TqHS8LrwbQvuHoy0h+U0v94Xlz5UckRsqMKKvN4wuM1sTZ3g6CEN7m0bsT3Dvi
muMczq8RUmR3cOGjJn8eL5KMJjye2B3KA6VDShE1oaPB04ATQJf1AkTK83675u3R
BA/Pu0erMvKOSABKIFmwjeRYD9aKeoN/lv7zdu5HzWWGTc7QV3SO4L591HRNSb15
FieC+I5tP0C9eBhJzZxUBOKTqIVsHRMzb5kL55KfNLvd1JnBlAH4SUa8XxaGLr6Y
62P6ruIdqqEsDITvKScgPZLRi7IF8nj3/qVdJY4UPA/r/9hmP4wwNrYlQZ02xCI9
NSLH4hpF+Yfj3XqRJzWqwVlWTPTo5VaTL9bGlqCyojh6VfhHx46pcX5EExvoJqaB
tmAHvjko9FFTiTP8ZaXMRxaNmyUgNc7K06WEbcs7G8dFmKUA351v0r23dlXhqDyS
fqNW/87x++Yy1SrAdBVlgl/Z5zkpu0MhXyE1pA8fs9oE9OWuO+OmB9lxZAO1cXkv
WeBpRpoczBJSBTMYW6jlf8B6jJznzIeDb3SxIOYCZv0DzSw2V7r7JkchNA3OmqEb
qDK1qyXNMUFtFSY9NuS8gmy0Hr8u6sTMxauQw4rpZD2ewMihAQtpXVO6EXS52XsT
65/ooLxlCm0UhZ9upMaCNsOvJs/PMW05mqX2c5DY6G9rIPxIs82DBlzkGdAjThLK
LCmXMfRg0V2W863wvJEDtXfmK9PT+oe9KtQX35JR2d2PwGdhh4GobhWaaD7+vn0r
geK/Zhal2+qmHwaBmMpR+UA3WSbM6qQ+PN0vIsR7tIDrLBoelw8v40dumXo/I3Z7
kPthLYg2eQ3tJLERrtnQR18oUdlKTqJ1wWOZ7Y4dy1XDAChd3140QW1yzJoFYfkl
8v4JKSp5LI8SqmgVhskeamyaBy8TUQSyDoHWBDSuexyN5MHOjVCSe83/alKQbYJM
nqbR9JipQTxy71AZkAMlveFu+ae15+wzzEu6vIxc4dpbMcXwHh9g4EU1YpNeyw16
t1tlrqzPJVCH6FZwu/Avv+i6pkPfvvhO0vSBy0PtGz4AeKyI8uYlhbrQCV9z26kD
6PP5YXRtHR4BObWBwDoDVoskDixlbzcP2grfAQR9vxfiDYtoR7USArK9XmjKZo+F
6gG+Y5cRQBzJYjPaoFOq26zYkMEUY6gDVgFT+9LFGOHihvBI0XILQEVQ6w4QbyUb
tHTYKvsCqwrr4BO/qMpa/+Gu8fxU0WAhx62QEL74JENHX8BHqHkTOFd+S3taysEp
o4wQJ2zBn5gUO2kySY6ugpeMYo86i4MsoXUnLO2vEAI8avaLmWMJXztZEuE1cEVn
Q70fTxHT/pB7cGppCYjlnZe6iB1Jdlqk7FayTutd41NT0ojM5k1cxs8+Z63QEZGL
dxtj+K3qUaWwVxcrcM0DkI0YHGiOcUZ7N2v7mrII/YZphoB7+pLwr3R3WMh+g/yr
qgo/UY/LVXn16h3RJQ7UaLhJ9baif180tVZB1C/bDCJPqCg+5+k/42ZHTXQYJnWY
z0DxI3my0qlxNB89smNAfBYRUEO9HtOCgfn/DPHoLC5NaMDDbIZQtGWJMwSD4bv/
Y/iC+zyISjF0ittjmOTJk6rz4JGEMzyXdKKGUuhjq3c/BewFkYw1dyAidTHgHEDN
GJL41b+1nJ9dqEk1ajlDF9mTcbuwwggL6yubKNeItItlgJSPF9ZHr7sSsDtgcCO5
Wo2dLbzmNt3QkpnrD5WXgQVb2GPt2guZM2FFnr1F5rK4ziu740S5RDcLm8hWLa9y
RMX8GZ96GeUKZWJM/lbLE7ykfWUTqam4sRhdnm4m5lzP2Y/6ptNpRIKJ3X7dkD3A
GDgDl8YkKUk7FBXRThuA6xhFbO7KTQjtYfhu2TOROPfNddznRAtM5JLPPDqFqV6Q
kvgAihK0mN0JLyrk4ATqmSa66OLo1krxINTVAS3NDwcvdLhOB+09wYYCQXYgarGQ
IKDH/mNzny1OJEa/1bDEWsXh03K35KoAy74FoxIvS7WseR/KxcqRenQf8lLpN8p0
6+nRtFme4H2CH1McUzSPVrpiBxSbI+LmpV6AGFJ/SIxRfzgyqA3X6ZF0VSeMcMer
S+viyo4aJYZvWfzItz8z9dKd9zg5D5JjQoUZQWIo3ZU5BNBqgLBalX8WQh3slDuK
yf8wVAgUERcYFxwmBaJRbMfVIX9HPGk1Skdeojazl94GY9V37RVMQ/IWxYgxplZi
THhA+xHZirsRGjgWtVBe9gp94ZiZSk9VQIIEiJiRMUTYC2ALQThiZYhs60lcOtZh
q1t0sjOS5pqVLv0q9BcX6gpXR4Fb//vloVRG3ax4nyba60gA05HV1yTOz4sJXS3d
FA9YGru0iRWzv5ersPTL597QL6dM77bAm8Fx1Jszk+/xn3Q4TbuhMZC5Hscbqj5F
+7od54cvN5zvWvbcIuG+PCNup+Q3rDVE0pCm8qhQr1Uql/BSaie8xnhb6wGt/Ivn
FynXGuo6cAA7gk7u3TSI3AngeHF24znMWzyoomktf3SC/hs1ZcBns1u/Kac/79l0
6wMt5ugxqnoyDXfjy8AnVYWJo/ywF7DzVBP5XiiO//4f3d2xK3yXIdJ95m6gAaxE
RHueiLa8NeFSC89KRDr2Zt+IxDTEW88tn7q85CSyyA4iTX4DYubbGWIDnFOqY2vA
+Dqd5eT0E7DaHG9zuMagbLG8qH1pFL9J7DODxBcuPer7ImUaV+aALRyfZWv2kinm
uMKc2o5eGCRj7kDyqWqZi1fDM5UkVQqIwkRWzVsXaU2UTu93hS/zRI4EWMQ5SE14
samxzl/f43fk9A68kl/rdpAxVVfz56chrBNUSpXkNhzUA0Go5Y6QiC4zmE8WRDB3
3Ix+9NhH38ZOI2ycMineHaWDZjrPVlVk/3C1WqVYfXdRfc92YEaB3xGqhozoSC+s
fWzdbteUqAjru1qJcdBnPNPEBRjdxUWO6kgBjKIHV7oG+jTbqGXjCE8SPiuECkIH
EftYnj1kJAZmMwnkTQGCfSccFdjz43SLEExxbVK5yzPEsly+lzLA6aoy5GXA1IBL
oSbfhxPFTycN7FVEs8VKvXOHQk0/Fp55tXJMEt30M20fHAz0XJl7fDm/ie96mwUw
ClXamAIENyj3yjyo1CVpYeiPb20I7+QhY7gO7VmflY5pC/AF/qqievO9Nslbdd9R
nUcCvtuxg0ywEjmo9sawp8TgrfiqZynQAJSiH1z4iSd8AJL7szzo0qP6PsRvYV7o
5TQMA7PftuStosKQz8Ew915z5/RgS0d7Sxdd/cAIuIw/lYxGpISD0aX9zEzxMWer
btwxu/saxsoG6GtiR1sWkWHxBTV3wHkZcPE3bHio435Nt3RY10XsfgbHmw3j7/Pm
YaJUvhFlzNaLBwi0nnLhljDBFdW6xMLtOnXrdOnmpw5egq1/WwOwEqIWGYvBRaFm
lPt9wkqgheIHb5UjVLphdwuA9u/yJtLjXRc/BQqjKhD1icKIrisHqWxj/SsPmavu
6uInQPAWP0shgztkhNdXGlP80UeenaNcr3FNn1cj3oDMAnUMuXTiptBUBmwRUqns
oLwcMpaKMn1gxx6RqoSt7iNOseC+PI1Hf06OiGbYcdnpp266aJL0txZZ3Ha9pwpF
0n35aYKWqBmR180H0xaqZ7aH0OW+jBKYbYremwq1KWNHHEgPTy0IQETMt8MQj8bq
SOZLuG38jgCACyr1mGTQwxiUr+3RrdCxvqLzXsoZ6KMxacKGH3WmawJGyR5h16+K
gzJ4GMWBF3KgAOiV781MgkQQCaI9uFvr/DJLoSC5NIrtie1vqwxMF8pmrtabzmNx
4zjML8I7O0TGHQa7sKbjmFsvagi/sSKt9/ruvS6CnoZbfENAwaM1ucn9aGq3qm/p
FBv3FIRfKmFnLQvCkLiria1bHpE15noMRgaqahg3cwLYt6DiF08/Ka8P1UyiwDoK
tNpOLi5nuFSuOtBAkQBDtgoJzAuHe4OinqlwSIHvA9vgZjdVQVIEKKMTdsmjkPRl
FZyGujSsHeac6AE2Ds4tnlE753VM7+pNA/1lSZNZZnmuok10Sod9b42irbKyEjZb
kmiUQ2MnylvN9qN5j7KoQhv203ivd7MWF+gVuiUWchLxWUPQRp7y0ilq3NjOp3HS
XpRs3PFUROiOMDut85I8tO/4aINA8uKClokOzD5P8SFeFHRZwaIQgS8yQEaoalNI
Cktm37mCR8TaMEX2wBIdcdy3A8S+rtnYrjhgp0hAaExK4fniukzhsrkJwPNyhISe
jVScRH1wjGy3Bxkq0o20bS/bPh+SRu+DytEKlHbRcFOd1eIDJi+BtWsy+ZS6DEid
0jHmytmafROumqxYcuG5PkR5/4TxFjbMUhxvAqN5JBLju9gyfrKxBMOSdRREzyAe
trCmAIeqOlW4zikwgqDxEY1p2SXcI30Wgg5QpDoRrr6uvpICiTXQ5h8h4m3C+a65
kR3ebmX2Sg6KyHL1DifJnOKZTANwpTpmpUIeuctCxBmTobABlAYeXbAikUpb2qja
rBay8qwl5tb2vB/beoGqZcELjnurE1nY5LQtcQ/eZckB+WhgXkFKe7yvzt3ZO2tp
gYapc9wNS2RcKzgDf8BDUFUaX7dbkciDiV+lacDwSQdj6FD5y7TiBYEM1wlBpqJH
lm8R14r5v9GndHtcV7CaqOM4Y+zbAejWlCg+Ts1ngn3vjcy992Ho85JKnza8eUpp
HDW7KN+dqbnhZXZ/K6qpXuoampx/cI8MH0igEGoXRZ/umcqVN3kzTP8UZcktMGxR
kd+CeiZCUZgK7yOu6q73VlbEBVPn857OJ08/RSVzMGSu/t9uZm3lnxCLpV0/xFIL
rd9ZgbZNMUH+6x/6OsUUFIyRWAFbm82N1BncQoqNfOGGIIp4xMJag8VGLtKiOvsr
lDNUKpwjLPZs37s52mUdcEbnm12+E8KHm2quvUN+OYJlRt1ZM9/dVZKMzqf4zJpu
R/vbFIyTQw8K5Q5haIAcKufSp80Stv48X+TBM5ePP9ZW++jNFK9h8E+oBwHiK6n5
00LuB089Sl4XIoJgczHnztZXxN+rnBmeHBKm7+WDrATR6LrJWxVIRaZE0QCeF+XC
siIBo9DhpSzX+YqksOR494AR6vhXQzv7lWzgLsPYnfT3O1Ge4rVuQeruUV8z5YPr
5V3qNTrAiLX2NbheJi44U5StU3VTh379aZL0lPo9c6GfZKapGDoyeyafYnkTODnI
1FSHXdKxVnMceuLtKO+NkyPZAh+atxVfrPaXlAunLr2uFoPRG0ge8i53KWx9jA1p
KGbhC/vqdSC0LNuVd4tTM3z2am6oLhG9ZSTUdT6OBbPCKgSy3eWtoMg7pvQyA/Ov
7VdHXnMBuK3YwsdBtQdKUmPUt/FjLbJs2FnYIMujz007vJ6mBFxRmzEg1bIkdF0x
j33whQt6YfOOzoS+Sg5AQ8jvcX26c5iLd/t4lw11m5jQforULUzLoUbRib/H3moN
zNtCyheb311DqYUUzpK0G4N8W9wvk/6jQT9MoDu9LczL9x2tSO2RhX6yN6mxHnW+
9wS1t3/x/3GwB8mFEBxRVpPY63eGcCwpJEk/Tp4JReS5GTrbORY6Tb8RU5g96MuF
yLyFqB9BZDJbjODPP38ZvERkKaymY1wNYEFTeG6BpyoJEBfLyqpYjC3yV7nikrr4
qp4odQKUVaXs25ec/lUfHyG23F7Zcwnd3myY29en68bM5ysYwK8AY1AX4XeYMj/9
3qBYQTl+LKG+lIn3Yc9sUggE4NZ/GykazKXqIdQlzxDEgGlY3h6NLKENmoENNxBt
TwTTVSxyASLTgloCt7sjdSoyK1q0kKLeFlNxqQPe9kLW8uqjbjDj2axN5AKxq8Ev
VvUGvhzdGK8LzHSEDREQafNp6XEuyXiNhjnTxU5JTl+pyr8QoIInKyX42y9diOu8
Nu47C7d7zQMa3ykpIVLhoNREm4GKinwCew4CgnpuxrNqtp1/uqHydZVWmG321AlB
1p389IsNsIsM7WULlWCfptGzI5+6OOsMG8n3CjJUVbDoMvYw+ecs+g/Nkx4//5qu
f74Dv1NenJIONCJHQBPSNbbISLuTKRHlXThEneozi45+fESKPu5gR400safGRvkN
NfkauaDwKWtXX0hwWqT0y70/KObmk/pvWrpLoXmlYSU3eksoqEYrBIxcT3mthviE
OU1Bz5eeYNFK3wm6bjUZwsfE8IUPIEanqNxyB7DOFHBiov1VzZi2HBBcMqbFZJnU
CMBhNKpp086hxsKkB+lJSJGhrqwmh6wR3WlbI3RxannuWCsmlEK+Gs9PUu2YzMQE
8N5aaJDftzuLisd+USuB7mzEpky5/VZU/jLnzYCY82YvgZgHXFOWJlAvr5V0I9Rx
hMnlXpTfBhSllZMOGlwAkgCCsYSzxIlLtHmNnyzzUh6Ry/JOxdVO0o9TOUYPYsPq
Vc7fQqftWoRDlVDkC0OAjW9G0DZf5JkhcDqBr7cWRJov67YRsL9uY1SSBvFjFv8j
K6QJOCYvcynx2Zxrc5cOv1SGnlC8pJfIlBbn8+AXZSkQh3+TKct8go68/cHMl0ad
mhaPkJ0x+sPxjwIO6CKRdrNah+KBPongrWoeDEgIDNfjvGzku+HIuTXm3zm9PZbQ
D2up7KDX2ImKKBKNS+031TjZtNn6hjIvURLDSDw9V48oKIi0jpgEpo9UCbjldvEV
Vw2VeIxeMFJF/zXliceLO4nvI3Te5+VQmCp1zcrHb9qv7xJVu/aGPeHw2r/AJNQR
nnWzx/aQjvqDhMRIABDK203S87D+Uj4CFHnBgJczgvBG8JCsLW9EVWC1IHuUhO8p
CjY9dSSr/J+7YfUTfcUSFYDHTtLim8oTikeClvF1LMZe/UhWYLSKLFU6sftFEGgC
b6U7GIoMuh0IlyEz7vJCyR1zDtuKx/FpkMd6IsavCKkFF3MWpBNdmCuhp/Sr6Hyk
s/ADuF4/0Rzw6nlzOMxPXqqljx8pXQ9uUJpYmwoIsFyNnMiFYHnw0RlHYlVSMH7S
xld9pi+x+jZUnXUX1JRr0L2CE9hEzCHNL3V1ALa5rwwA8e/2j2EUBFG25D3NCOGu
fhQvshtKBq1V7em8ioPyxiUElfXSXoSLQ5KUyY62l9cqbdJ/arMycPaS4otSHct+
MFrM1dsCrJ/mWDawYxeLD0niSVwIG64qjNj5ZqP6OZkJFfjAQKxMIg/q0Ce0KDH6
KUoaP0n6x8rv2eNz1/vknFPWmMKidvja/z0jAUE5c9/jm+4B21rDWcBzQ2DastHm
PocjEymxYxWiXOy7hHkJIE+crxcv9DL5ippxIB1rOifRt2YXlz6PXAtgGZ0BZ2we
dRx+CbLf6ccs2m7YPcfcbb473WnbvdiQBz28KkCeUI1wj7UIg1KvjWlT3rBhPzqm
rrQYyLwfzufKYrCvt4FMEpzNgJWo7Zsozft3CBNbZb5g1k7dzL7JsAwx5xNazzGZ
RuDqc+a5l3U7t3kxbvYpwssnEzqj9tpx/LZlt/L1+8oG5cfT5MZmiox57wX+e+9P
x1vNKynE5+n1R5YNsK63HLvFSRVioZl5J5Wq8ZUL/PYUvO4urBhTM3LMzRAW7ejE
lC9URKGs19b2rwJ0r47WyKeNd6wQoOEtWFG69o08hy5BdBvsJVfVXRtKPWyv1vJA
GLCGWIetrhVpf+h1PV2BsR0VHFHC4G5RP7Kj/ffO6xH7yYRALZs26yLGMAyP6eUY
65I0PengVB1sG6VH80+DqwxTa/sK4SOyjt1yQ2wUG292fD+owonSwHx+JS87AAX1
QHR4H6HtPlXEaoZuljuuYEDzkTYK2QC3S2nCp4rT5yCCTylEh1+aZbu8Vq6qVqTp
qPEnssLkfSZjpkICetZsowsRkTqxTTVvPr+xDHI4DZauo2cvAd1fd1QYWzA6oMU7
yXp/5Y4jWHdnXGKQuYh2IKQgn0foGJ96cV8mqJ29/EkyIXBIuKQB4M2C78HZK98y
9zpfwBATxaLrgmWtDNPB8ura3ISZ1jeC+ARPbW09ljEW4OgERmR614NopBY51GuK
IhmeML+303KPEm3inbjtbPop7tlPz1W/CJF0ZrpuSsuKxfbJlwDrd+lUgMzEHwTs
2O4F+pNbfmmS2N42OmjX3ly0v8ABE/FdmyGY/sHmh0KRRw08OCvTT4U1GRo2Riny
eLI5JdrOLr8fKGOwSj4FBp3RzDql1/+xiGmm6Bwk1noHgI3VHw4Jn4kvVcvmDzXJ
zZuVE2akSvFcgeKeqpGoAPg9cjfNhX3XZnnkloTNSmFCJa/4b4gf0sQJkhAkB9/l
vZIJJa6D0GqFrcdq+WXFr40chqX2zNuJNhyYQl27+6JjFN9Vm2MaCTnFuuPmWXRz
KSpwlIObXhuSf7+2xr+WYGaAKKUgi5PG+ddXpXT5PJTfe7sfnq3IqtQC2H+CEECF
OFPhUOaA/t0wyupdWb5Lqz+3QRPEj3YRiefaV/T1crJlURduuKuRIIfEE2zhdqDV
t076ejBKJad86O48L5B5NI+QXeGzJbedWC2ydyS99YiPYZNoH1YrLNNsN7sWMOoe
3QJH035u/+8/zvobFz7TDmCasu897nTc/GTz/lQUt52SJdUBavGsKpd9aQ5Kkp1N
vZLGtTZfa+17za2WvclaoB7/TT/8xnBJRp94lJbB9fJTIWPxdh7GjjCqZkCH5tH2
XSrN0Zo/9J2xkDqpQacGMhZowhxEx+foVg9c4S+g8xS94DvEKubfZO/BRlPY5gOh
k4JcYDyqh/crHZ5kyBdOhTEtpGRdAkN4xpEP7VOV98o71ziVlCHGnwzsIIHDR0F8
5bvWJ5oB5+YzDcJ1Iq+WUrywBFxvYx5+Oq3hf1i5B6H1bH/+ySgHeJZ5cd7wxTT2
f5OytQjCk9QTCerWlcINnwTIe/+UDcB9rFq4H/p8jv8Fl8Q0An2rtr8k9XIqNiBD
I7VLzH8VaovYcUV3uypX5H+9sg5zA2f1G9A1+eWDu4EJP+EgqdkPmgj+zV+djdGP
NnchBpkTeKTtASvJBZM130UnJNhNZa4ngUJK0Qpkt9lyB4c0q/UTDH40QsA13JbF
NEa6kyNVE7bcbzebe4AThKBRy+NZCj1Cn+WOvb3yByG4PAKAQPYpUfQA7Z7wTqFY
4eL5vU0wV4ArXCR7QKp7Y19CLv0FTQDwv+tr5QZCnejIbIHME3ADU48Qlgop/9OV
BoCiBwD9mzSRy88XwCALf/zllGDX5cvFNOL2wFZb+a2NVHwBXg426Ck83i7CvAjY
O7YNglKXb/gKJNq2c1fagG7ewSVO83GEd/rObQvYsW0eBUOOe7cQ5uhZyueLY8+d
2nOsiAhLu9YhokmI0VyKpKH4IP6BnMGz9MgT3fCFUTI5H8tQHMrvn+p8mViRrsW3
s54f1uFJt8XevyQBJrIFd9XOMv23SA/2ZJYaDIPp/eSXgq08SM3xyc7eJejqptmo
YUxyCsCs/xUrQMbcetjc09Ewdi+clNNVueuqBt/q4mC/3l9k5Blr/VAQsC3EQTUh
uaVZuqYfXmmbwtafswfRTjtpLxuyXuxuYTfG/2GLNLSepDtw8vnhHMKTD6NuRIma
hRunAGPCBvzKflF8FfPxWpV5IOLt4WVFupm7TaZWhrkQ5W7NUchM1drKm8yx5wId
HO1l8897ZTLp032hJhXkQ6G1DUjlQvtCP4FQNpN03QrXZH7oIfnDVxcQsBJc/g2s
6FSa3OIcQesum7mptEBxKDvKZhevqkokPQo7SbHeBHBBkg80SrzKwqRQk1VrpzZ7
+50hvKWs4dg/G+GtPOVkgnf53zZA3nuEC4BpPvnfBgi6SelH5t3JtMO3/Wq+ew6j
z4ym50NAIuwtiTz/o2riWmYevL/8OuyB3f/A6OtstzU1lwNvxk9ToMZ6MsCzjBrF
WQqh1viiJRZQ+wYiMsbLEYAnFyeF9g67otbQCrhDAYJb83FWdpojL9SUe4wca5zi
6yUtiy/7ZN77ozmwM1vt0eTJjUY2UpFG75jkaicXN4vrPTvwRJ7UIGzdtxq7e0Ec
K9D4m3fVbnFvs4enDZwt3I87HFPoxhidSuOmracoxu8ACY5MMpYFDHydLTZS0nNL
Uvu+kiKkes/mtLYAqF+E2VXWsa53lOiXU4PaGtAtRJ/xDBdKCgQsd1hr6uHfSQmp
rhPtM+HGcaCjRHzt2vTG3Xe9qdeJwR8twjm1kEgmHw+ATPebgO7q6Bncnpg80boI
APzeAe0FaL2UXjc1Hxw35r4+kRC5A2hTzuUhCjiFPB/QBZWS7/o7u+taQQKLYBuu
yEbN6m40KdtZKUwO3XguHm6Mu7088oDTaghgBt14enOJ1YA5Z9/vtkN4a+fO8nLX
ELyZ6yOcZvWnzn4g7VW5Oglu3RTj4E89EQGRdk5hZ4xZvfEs2t5emQ45D5+LgQt8
HBjw2CMrl3Zb66ADpi6Y+fwdmd+jGDoU1/vwRZfBnKdCt1vXchndVQx2bgRqaXzO
l6osaNVmXS0k79ZEM2HU9IQlqx6sTccmQKNBK9WKqS4PkobGyh3PMlTpJCMe3DZA
MJng6ijfOB+5P1YFWSqJksIFtUFEwAOJDsQCiNaSR6r4Jl0XPqE7JO+j77DIqHcR
FL0HOAoHBIjzh2Z0ROp8BJ/HYeJsZUzHGjuadR0CYPA39Ww6CEU/TV/Kl0g+aheQ
0lYp03CUIfSg9xw6TylkPvfGxLwqAwwPQHd8HjMUQt89Ws4ABhumWFsuErhvliiq
EVfjdfdeal3Ei7VvXHi9IO8RJsPmom8W0xFcYwl8ErynadMS43xegGDDVeLGx99T
jPHHEHoYYTTOC2nFy9/nvQiYrDY7gfpNb8Az3wDV/XjfCMDt6JwNFh9FMRRBapuU
xVZWPzdo4F+xeFxjE7XOaH7GSdC8JN/q7OraxR1wPfWdGd4EllQvOAUgHUHvQ5W0
InTRhwks+kWGuxY5dt3VM9Uo4e5SlFiAtsIFufVykjKY7LGM8q8Oihicf0lcZ799
Mt7ctAhq8b5tZGNnwQMCO/V59pFjm8rit01Br1Jp6OxUobnHrT/j+UHFaMSo28vj
8TlG9psgAuHie3IwTE+Bmpej2W4Y3glRqDYe1Zu0brQMscpk7C2G543nUxZCX8Sz
p2aQgwOCpZOUXZY4izhkNnamoWYApRsgihwuuKSNY/Hhh8JtLDgCJiORuYWxoUHh
Ao+eicjwGe1sYztQ1TSsnv0HITPhmBTSMH2J70vW5N+exnlBLbZ83GOcU9sWM19S
cWkqH3/Lq5G68R/FoQP8xqXAT0Jny4y+WwygwQm2JaR+99OopxheL42F6ZYp9lnb
cJ7WZA1zWMX8ClVA09v4Bm+co8p/VZLLZGo3HFWMOFRvXBGO35DX46tO5ighxkog
zIskBLAdD2H5PCoNt7pu8KTZnX53NIJbA+Y8sNTN2ixeRU9DXsrTfUJtbnp4yx/d
QPz/IJ0TaA521wUUM3pTuQzDOXycAE2v3jVxrfFlH3ilGixWmebueExQW+LFX1zy
5Ryr8Q93Jq9ZhPBJOq6hD3FqkJ5AnnFCZe7q9Mwa/BLklrwqCrRhsb/NnhABYNtY
AY0dmceaEC0PBPEnjoE319GXc+N9uzF6BShLqSWqPbBtCKKa4Yz5P7z1RFHs8Wka
rGyrI00wNm8WZBNx7kFdWCu4bq9O9uXksSeib6oA95pMYUu8HZ/9aG11JumqgqD6
I6y78dmVIWy8BUKlj57p2VU+P0gQrbpk+Abg5VgVLgWgtj6jr2U0r1Z0NPvxaWYl
Uzv5faka7ivuB42rBdbyfCCwHcLLkK0Ko8sBd4iz0Dr86o+jV/P+S5Af4rQq4oQq
npKs38Gr4g/OquA0gbfhaLJDTc3FuMCiM3N5UJZOlW4gL5K6ZcR89s/eCnT8VAvo
yblUHtOj46wu2piH+s33g394UjHL7uWopyq2JtfqA69wkwlnqh/miip26F5rPOFz
t3ubBfXrBo9Gea9ixCe8gLdqk+qPYsSE4fzCzpIdgLdD+HtSro2B20PDKEmBCVB1
CPH0qYDlI2QBNOmqf9WWOJQiK2tCFF9hvP4PhGvj3bT38ttKakHtwIP+90T34Lm5
o8LV6fo9G/k+6UmhvnaQ8POmxNamwhtODBhhRuilH8coNoxMsiclN+usonCyX++o
u9LO+bdVTTd8dBX4b+lVVG44WZrUZ/ZyBtTIL8sXBGxmQ4gEsvmlvMjIJ7mlHx8C
3Tqjqqbbj7udQk+aJSWGXWX5je6X6JY8UCa0AEkcQFz/MnX/Iz5w5MHPIGSU7TY1
lhunvvdz5skNxvvofPcWieSTW5ZEUCBqXsuypgmM2zXtT+sArYlT3ormIqmYZYYm
XbD5bnAcZtoAnXrpJ43jyL3oRTViVH01fKgEWEtmJxJY1E3CAq777cT0bNxNEvcD
igLE6I+xmqEzJ/dN6qnRpmreRMWhK86u3c5m6eZz4/SQwVV+v0ZKR24qorHdKj6I
nlr06H9+bcdOSaw+YFN8LKBcAU5sohVzRk7kx+6F6fPLg+uBCrKZmag2hAhgYXf3
d1FqkUBaYZSPvY//2EXloKTE1pUtH6mFWHuCu881J6+CBfmi1i91RMw1n9Yl2zcW
Jyh412UQlOFUrbfxVSjJ7V10idwodWkPSVwwpVIgWhz6tfckiONuB+mAY+9IHn3F
m6148Tzq4fdR99TzLvA9QevNB2w+HBEl1DBvt2qkgusLR9UCfjX8ngbaRsFZgDgP
eUK5UwXzRmFtfTdUBmTDna9Pi92UVLgIp9TCnag3FhuyxZ2irTSBRlvihch/3imx
hag0Ln5I/WaOZUuNqqaiMWJQQH6Gz8qvn0kZnRwNCK2Kl+Hrf4J1ICzyPXzAeYBp
qUW54S6a/YMMpj2jHnXEdWEgl8YJNydfh1Q/PNLIjRSKzx5w0sgRc+B61CrkTN3P
IzjlakTLWwoFsbLYbqDhiEV7vgepMcoK3v2b5sK0+ydL+ho0vm/IuNUhJUxucY47
bLGsWvS05bJxRAHX8C4BdBjoLZbOzx9PowNcZjM5DQ6ZXjVojGR/nG8Pt+UGcW/R
DYcH64ascVCOmlpUwxQIwTYqq874SGldCd5T/GV5thVXnTXi6UeUg3ewFcoex8Pi
9XPtvijYtiF1L2fVQdyKfO3Q13clHpIpJjz6iJKSg1oGx/zzO26we3sJvL38uzKr
WWvmlNzVDjjSKxR5piceRYj4STEvtcy3YNw/7N1yVtLHoCqtBqgo+FY95jqwCmAW
pG+x9XL8ifMSmzT1J12PRzCanfsD8ThqOZDHYahlIBvJIF6Bkiv3otXutW1baEZ0
TZc1667fqaa2h0PP7WusJY+uiQZHtahuMa0pOQwXn1qcyMRIEkDS73fhmVKN2XRs
6bxKaqSdOQcLjig9VvfDOzY4IPbQcXRE+syfscJ/KKnMDFwgO34/VIl6Bi1vObfj
A3a0JpeuDsgIRy8fp4VwGudqQfjDeauS8TWY+HmFaBuv7RPAcJtKK6hRhxeDl+4f
8hB/o1ZWn1pdJRKzIX2osycMMaerZvvXoKXlBiP25nB80kgDzy+4p+0yawouHQj3
O73LmhWHv0BqS5whcJSDHTVSDr4vZBaFWGrtvEJTm3YBgp21PGhEmv1eGWhdmGUf
4lA760/m5wmlT1EzzHlBJVP+BKh6DCwmJh2RxtdPrTgLRL7oyrZL116AJvfYigE9
dBpY48n4Hz01iah14QjUatbzMm4KhK826mxhv2TeAFgivvZbz5CKS2K13+v8iY2b
fEWQ9LhllBHc9lQheqIVAFG8UoLYnfbzj4oaK7QHZkLc4G5CH2MafBP941oSGvS4
IZQ0h0iNts1DVfhR1octlIbqySqiDhSNzj5iSjJJUYPCoWS/ahIVuhOtYGKgnFB3
6O02uFCQOwf9Nyq1oCX/VAgMwBNWpwflDjOUEeqrFx+ZW8hsgFpxHn4ysluWyy3q
3gBr5fGH2LfVLSywvLuR/sA/a9lINTh1FJ15nKL8K2oNdxmutHtucZ4UPn4G7Mra
mr8ossKDkJRzKzjXJMD90TXT/uBd9Fhgs8fRlsOm3lquZK83cwvsXS+qljqDnSg0
cA/TAJ8p/yJFMbZiq9qmZWGTUynzif9NUJ4mR/orVlf2AeT/vRJwe3Nz0IaKKtYl
io8ge1SfiQssEJcClm/GuBCgRaW36nqJmQl9D+r7VGsIwt6HgtopitcY6L8Vt/SU
fvzxux39h7pnV15xAxoVwjm6wtKSrG8NgaeQ+et22tuZKYuMvFco92A07eDbVCA2
xqPDIk8eWykCJdaIJ04tTTEy5kuEWP4uQIGU+lNxy87NPlrAot2snRbWAw7aG9PC
9dljbAhBXqG3G0aEO0/d8hf/AxYrcg499dUGU++lqpr1KriB1Ihb0dhEBerhTmFg
1CbfH9C8A5QWg7ibwRCDHDZwd/Z8syoHWqayElG7fDEzwHGbQpuUARhnNoNZ5dRO
G7on0q6DW0mTg7liw6bg1vdIiKjUtle3Zs38B8cI9DClb9Ny0tQHXTQVY9Fgs+6h
K9tHKjdfWElLnlOO04aObb07DqgoSiRxcODfNxEDQDOqz4uuC4BWLB1k1NwcI0iN
ESOYRqMa1yVgoNqaet/l1d4qRjk1G1J2yUEsFWR+6fMej8yhEe9bhgFDTLgjseW4
/sy4i7QUONElzpGvM22N1M3zTH0IcOo1DqOHZgc/GxatI9kgGO6Hdy025TRxgEQI
3CX+tlqGwn+OggLCoLCZliZEli1n9Zso2OasXmmiQEGdgMpTM5nz3UuHeQqXRUp4
ArE9gj4EzuW/HUB6zmB8rvvl/Zgs1Ky62dWqFQhDb9AumWfr+1FCniVQK4K1iZnu
SCTJQnOnKprfE5w1CVBvKVOhXtf88nCjkKMByZjwn7LzAbiLL74e/OFC1BtqJELy
hkhygvDtcw1IJJTR5sYEd5JjASkBlrY+sTjkyr4lHln2zZ8iRIaYwhgLHK3/9g9u
q5JwGJnOLwCSwjf1et4gCKuRrwowc/2XywuvX/pkY9LUZH1dtGESVbODZ11FOhvO
nSiJJ+bsyhWDEO9moWMJssaiGmkufGTzQveyLWILGvtYfYveoTaCubYxKx1/I8lT
jf5/UETQxJOCn8Muv0VgS3bSfVFRaK4jYYOxLq6gyS4yLG6XPgfS16UIIchRK8QR
`pragma protect end_protected
